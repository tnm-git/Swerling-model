`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2015"
`protect key_keyowner = "Cadence Design Systems.", key_keyname = "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
NTHUp4mVkg7HTDVRaDSCHpzyiGedBWFNYCLwSIF/r/+39SCtPkOkLMHnaz31+3NjlFSsUDvSpZ2p
DZZqZOGJEw==

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
Ws38mdxpYlFdBlEevfRHjWoke1gjCxGPiM4B1lJwmHi3XfZKznin3sI0Wb8K6zkQMAN2ESHTtytY
sUCZlqH8J57dUhzKw0buc68LVgXFC9+PINzpRLT8UJJHeWBh7JdgfFwNYgaRaiPJwTebwAAdiKmf
0ptAG3PntKrBAMXPXAI=

`protect key_keyowner = "Synopsys", key_keyname = "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
Ofbv0Kr/xD5rXpVONXsPFKph9CYFvK2F+qQmUrkH23twvmj9MT2E4VlUlEW7DR3qHWclOzR2zdGz
fS/5JUHaIyPRFiIACQusqKcZlUr9aOFLYLZEArg+cRAYul9ShRppwxxLEyR71UGvWZCQ2Z/CIH3A
+odZjekmbujgEQeMKdQ=

`protect key_keyowner = "Aldec", key_keyname = "ALDEC15_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
M7LPcpqpLKsYYWD+CEkS5irzuJpgpmpSyueYxRu49wliC39VnRZ4557j1e6+oJw78WZ/aznyCn2U
J08/IwSiO1XXEJYf8HNaRZ0uu09spn5qOqzK2FslQMimohIbyTt/CdjNaEh6GFQyORcJ4+Za2TLY
2g8FsYYfWar9JvfI+XXj+dmmIOPvNrJ/qzelAMPpSmg76MwH8V6JVClgh+zbLN5UMpGy2kGxwtIm
EALWX5C/QpOX7i58jcjhXdWmZJ2i1fL84rOk6YWLsG/pX+oGh1Z8JryE0XgFJqabKugFB42vjsW7
1zZ2gf1bIYpK9izin1sO3+EUU5vVON3qKvUHsQ==

`protect key_keyowner = "ATRENTA", key_keyname = "ATR-SG-2015-RSA-3", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
glrJvcXyzp2EzL/CLILnzfOrTLJ5SQ/UQNv1rAy7YFhodMmtlkAjNUABFZZbCUYKZB6Rhl1udnEw
21Kv698jQrb61GN+C6MamSzTmRu8AxeXCbfJOE0ABEGL0tVv8xCeEEZYiAWbVydV5oFeQ0aUx0zO
dKIjvqNzwHWexe+YZ+P3zcHwU4tuJ/ZDiT7cQeOwDO/OnDydlzUxB62Grp23yRbR5IPKsZnzeEky
LQaxLIdNZ/X1xNacnSIcyZ7CssjWZkX8eTteJQ8/ugnmlCMPLFleg+erqI8FMELaNgfsdXOhmGHb
1DgtGFVNZrSqpMUDkq6mn5vK8lXdJMtvQnP8QA==

`protect key_keyowner = "Xilinx", key_keyname = "xilinx_2016_05", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
UNY4I3doME08ZZhQFl0GsQW+KS3EpG5s9WXIBDDgt4eNqLeTR8m404YWwnDjB5GVUe0L45QTW7aE
GYDchzaVHAt42l1k7dU93WpNQI2HYFOu/zbUNyg7Q60rmMVIwMuOjeACc8mMFPlX2F07Ao/qsre9
7WcMwYLHyYdn+XVyrTtwcwfLADI6E/lLTMXYnZm1QZy2wz71Irf14LQ+02Uz8Cknw2PdGF+hwrvP
z7giPbt2zqLNA8/+Ht3bmEQ/SDHzLIPNyNQ3cIGffVu1RZv1dkrTFYdt5icKcepEDwvUqYhUvlPt
zPYpXsRhh5G/ABEWRJnscmXNjKGgKmc1mvm2zg==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 432720)
`protect data_block
LCcO08qvaRfA12qrgvHpaQOsAEy5se6wPgtYra4e7ozmwBUqdaH0HeBxNlGIa/PkEIZlnxh17rnJ
RjIyqg/OIgkaIGhueH10/4rYWF0P+w/qArhkkVVPH2rJTDyjDez7LECB6G7FhJKekYr8iol5oL6d
U3SuTH4lSTXZ7vPjR6jM9Rsexa5cWDubwqkIEnzaINrkjx7LfAmTBEVhSHUVA/pYtFmK/CH05xhm
mMFIEp69XUE/3bGGU42S75pTUYNWpiSTxjpNHbT/BIgxlTJFZ1sMFSfFjQ9HdeUaQ7jbbtit4A+L
6/LWbZqrzkHaiHXKjyfvlfKtzsLFZy6bvfxfikeOrWpkBfJIPchjgvmAB0y14DHohPOwDXKuXbob
wpjXZ5eWQiTSGrXQtezt5wpcyDvG8NshFuQryC8sf8KIFb5CiQPgml+Ecv+e8Coz4wtr/xGzX+QO
A75Z7Bzm8ZnR/AiRG8h5Ttc7wG5fEGdgd1HvrvOp5PqvMBk9OxqqK4tOOQr2ine+zDybtuq6fGfh
1JHOaWphZnJQS7IWt4RiRJ7uTqshszHH344V9AmGe/SHH34Fr/SKZNm2Z+6AJzdSD/p1gSirMSQr
+TM6l3hZJ9vJlCCkXaONKXh0ymanPenO1EtlBsh1k3XtmJN1OaZDMZBUut7+kgUIiHOYFQGrI6Yh
treWm7k8YBxvw9KX9AqoP8YyMnVsmH1daEVGmzkEuDe5eynhkVHnYFWv7hNKYSNiYvyhYoeVfwzv
vUq8oIplAuLQ15hC3iWA6uC+7dHYtQkyWJimh3DGdp4PLWpl9xorDjiBD5lCzIcBL2ighAgX06rL
xwT0TwQZCmmIKKnN48ZS1m42HI0DByvISL3DjBF8rIaSokv4pSHVOxnmH+STmgt1x0o7f7lbtKZC
jA684/XhhKS1QJWcuC1RT7dKNxoSRK1a/fPC4E6/VRVSGmSilgY3U9xzwJFsMh02LBkJkMXrA32Z
1apOqG+C3+pAsU3MGS26YrCCc8BywgAjPNTcS5Xpf6R7B30ohbBpOWcZOenr/ZS46/UeQ4j9NKPp
KQisOxVOTnscESmpgBXdSJkzdoaMGruMVvhKRrEZ00nWaBlcDS3mf7Tgrvv+1jzxu2day2lSFxMs
xVjCwnsS5CngQs4sHYwey7aJa3QhSeY5OYGFPhLE7qhdvE3qWDV88csey70mfEa8a2wisQAfT2Z8
2ZACWy3DgErZ3p3yzxJUxHSBj3RNNbkg/E76HdEV0OD0J1/QuctHoFed5q3+HCXXc3vl0/uzyFRv
CSdC1ncC6R8QOJy1nNXJAzXLO0X0Va1f+DdJyg57uBw95V/xth13/8wYZUBUuBR+5VfpeJSY13Bl
EtHLhHikzM3bXeAarossDMA3MWQhVMkyETvRpkFJz6hwU+zIislXaVAmp5O/enmi8bcYJgu/lfOi
lERfsWvD1q5IIk678EPLAhe3Ge29oOSGkgAscTce+7w5f6eoq7RJuDA1xiyyHu3KYxCTR0hzf7tL
5l9tW31Ys+/wiqIu5AIi/K/UIopLlg17J+8WpRATufNNlNIevuIgjsNsz5dujeZVJ4C11wDSuVGH
AI1WS8+uQS2xljHiz4UfmItS3a4BlAxOSZKCtYEjyW0FIO1zR5k6eFUZamwfFbxUDDhoJAaQIOeu
MM5X/p6YqNfx8qtPUlpSv4mmXsiAI6op9Ww6ocXU95ymvWokQXPoDH9Q1mtC+vbGp51k+jmsOILI
fjZ1pQw+X3KH3HbnEPtrwXHteC7Cng9QI6cjLdvRleBqbof/Wybn8uGPLyYTHdxy0k6KXZzV+Yc5
eOl4C0GywrNBC3PomEsrPieauVv8gRAmxlAh2+6pvFkbWZlMvIlEVhqEkk1/pjjoyazzxOzEBH7x
SGo9xGjbr6RZQJVHAZZ472jiK2BiyKnlfwruuwB7eW34kLHtcUAy4+xfFSJkdcPXJaWXP0GLAtDr
2DJoa1qDOUAjmsG15Z/fzxn9l4OeY4pr8AOtNVFHpPgXm62BHdWPvOaQge0dwm7kTvT3wfNhM030
BdieWsXUXlqZs21W/CdmqhDpVjQwWDmxuqLcgc3xyhZsP2iYaq3BW0VkV4U342C7mqf31FMaIzxZ
fgjOracxdb72JVz2Xdj670Z0FYSkDs09gfSAfEPlgh/3naLULJ2tdYZKK/4PvbXH0YI6wvD8vzMH
SgivcDiK4RNnPvwOcqkuI3Ts6jfyDDpFFHbO3WOyN0B6IXsthmE6BTE2qhk9tZYD5WDrAEwheHmS
/gpTbtXMH301f2ymsBFocWz0nA2R30TwQtwbsoK8fKpV9t6dCsDXczHUBHM3ULGvXvXU4g3xjqYI
EpyCU6ggHLqvFmUZzVJXn4cQPOe6wjU0nybFJbrn2JOQ5Alsg3+BFcmxnfjyx0PBg2IRAIHOLFaJ
MxQeKEA7DngDin76+v101tLNiEqivC2Mo0/Nz9zXxek2u7s4O5jiWHdIaXuCd/7gozieUKPG3DKN
LJOd/5MSyHz5jvZSt8WzBg0r4MWJgVFYbJjhGDaAYmhBSWf3zQJqcjeZlI3CvGI+XXKZv7aOKS+Y
/LdomuCuPhrBTFUrfRf7YooS5oitc1xJE4qMImeIFLrlylo+ij8WaKtW/3mOgLLMncqa91S4+z/3
sdiMS5uQ4WA92F7LoQg1CeMOoNNVp03Fb6DABLUmQxZ+iKKV9mPH5IfmMX2jt8XcFyvSTUV1iyOh
zjbUl7bLX3pdqh9wIm1TUpaxCiBp4qTQvt1s0Octo6PGrj+UslCXw3XFVpinTZv/y/5wPLfeJ/rI
5YFp9vqRqNn5opQ97SxXECK4UtxuT58XgsDKJiLFbaOENCZ1vMg2wKMCV9jC47iFH4/aF6jC/Kqt
ZRKmBu0btkdU96ksgwsuQ+j+fUKc2loOdtXQPyFpavdPdLifqYDjtVp/ZfA4Vz32MdZKlmYgPAf+
OYSN7fQC3KwBksWYyBeSvkYgW61Rflvkt2Fivvf2Jdf5DZ5hxLURQQh/2X7vWhK/14flZr+Ipz7z
NHRQNT64Q4jv5eNf/4d3D2MCMKiPJmM/B3770AQIvr4JVHY8EE5wHloJlPy8YEiOHTurr6E6EUQ6
Cnu8UwCAyPm7DTLJ1MINOBwFSc0WQMUHiOWfrU/Xk6M8c7bm1ODSU0OsWfDiFxI2yKXEfekyZVPE
AaE/ugmVCaUyzsq70jqb8vEDzLAGkx5kHjHTGWjKDSXhaJpqUn6UjCm+gWpR3SxoruziiH8oYubb
k4n4m9cwCM7MNLuBQwHlsgpg0Dp16ZNuP7KWoa1JElESCR1wuQx79YuEc2CIq2i+s8I2MOJ11/V8
HKCRNjly0YAxvH1/MmrBNhqwXxib2/YyaMzgYNKAPUqp9yM8SSCfFvF2P6WcUpsZEvJ2X0x6X73R
1mSGSAVdQS2s3QJzJ0T62r2aehE4TZa7iUpIdg/h5Ukwhuq6uLuswGVEpOR64hrrb+DBGCCknoDN
CRmcBpIsPRX0PDGL0BzhX6gZOv0eBc2iV5YtLJxhPPUGjXlHqhr/XgjkEcV/q1xD5npkiUTQI7CO
UgR5EitA9GNZk6ZqJTO4LkLGsKB5GvImEAbS9I0GsNkgol4D/M2MrqsyWnPGtX+QwCJY0OUcjjBW
Wd/bu+GImn1ymFkNgynB1K8bOvwOAk5pDFStvIvln8CjXVGnsf3p9X3y+R7zCi2CyYCXclXKvMMK
RmSvMmHPbpVtj9uXnqxqrdKp7dCXVdojwyj305d4N3IfR7mltdpUSbCyQ3Zi+GCEntmz93+LiT9Q
mNcnR24jQM91fnnKgzidIkTlgTRj1mlZ6See5SlonzRXaAwS/9ZA/wf8xo6plirjwC+dsMw01KM1
J5MQnYKIOv4iB8ifCt0E9DBQv2s4HDtv1Jc6xxHHshUWAotA6HG/sNQHNRHvuT2JBsc0wugnOqRH
+mL3l4iXR4gU9Marfn5pH6aC23RrE1Hp3HFm5FZKyNaB0XvYYjDk+q7LnDbGIvqe3OlAjwY8wc66
02x/P/o9rZ+zgZdIBjR24bZsgAvHi8/yjFWN5g0isYcIJhd6tqah8gJn7BBvsiswz4m9JRq5i93w
CVAfmLV5c/8pUq04cjXjdq0B+qlmjFbF3Km27DcYJkQl1TWFFLWSjIsAVkn/cDF7GqjVRynTkGCA
4rMLEEtVeiocYfBa3ylrl8xJBfPy0YEy9R4jGSznSsQbE6YX/iBEMtcst8zRfifHV74wcAplOLSq
FC4NGqb3SizhhCEq/T1rb8IXV2pfb0hgqjk3HjjEd4UL/YbFZ12NrBaMAbKQo/j0DjBJeWEMDeXP
t2IBHRN5kYnLMsvCtdvwi1Hg3wOYyOYAI0q9GUzzkarlSQqvB+Lmn8cHWRgwh7t3VXBzA7bZRkfA
two/76BsmTaKYzX4hvYgcDUyZLhDgi+5I9dyGFy7CeQTryueoIAJ3lMqtQlLIyGspUq6JQkSfbAs
o0KUbbocHg4Ml1YbudoKr1f/cwyqD2NdR7kp5cH6lUDTE3Ms0qbWNyZFtifPasx7CEyAowBSq9gJ
ODEnHh1RaDOo5WWXwXBzZyXqq2N7G5V/AEYageZqy6W57oAFE3/k2cvJy/IhXMzbTcGGyM+OpFUZ
6PMoEUVtzochisBYaRQ8lRQRltd8l2m+JsjlCKyQvLPSznYm2FzwYxPl2S4HBy9/XvMYBhioaGrn
q9gxYrUytbwqr5jZf1+4T3JiRJTDYIa66Cb3Z5xIzeKsHf1vJDkiHQsAGKrYGi8MfI8GX7/IkWEp
117/t+xMjUsU89iROggEmzit8vb+ixzZw3Nx+wtDpNRCAiKjk5tQsrJKEplpHDUF6ws4svqW/8Y2
Yy8MCNSKe3YxkYW1wBOcbuKUeY/vVn6yqn6oNmrhNNlky5yF+nYrSaHEmCUWwGR/bAZlStsyVsZ5
s9tGvk1JeR8hMHFbSisBe42nh/jh8WBPTyHYjapyFUxcGwl9oH5Ov1+++qjta1UL0h9OBarwcz9x
BSju89uEJcJJPFReb7QiAONzz84yrqtSH94tPxXCjO0g3CpExx3pskpwPKRqbpU0xs89jBszI8t0
CbKbRfz18h69j2iHQvbilPFAiv36WpLYfYLVCIcm8xZnmWXS2s0VqDAofNYkSzWKyS+bbRLMNCHb
y4GK//mYIyH2wnlCRYZiNEJVoY1YxCyWpL/3OvY8cYszBrX3urWqjg4SzTtKoXCYshnCzgwLsMDh
MwOuZawtmkH5aT6qbraH86IhJ67/aWVG5hDDKxM6OZusmntijAx8cit3LlW/2wgo3pRKJkSYZobi
Can772nrVmDLH4pPBT5fRwK5Bzt9mH97P+UM6NNOclO/1tygxxqCGK9mxHbrFZL6tNuqDay7xVEm
chWE5mBCxjhETjGQMyUTLhsrKWrH9AfA4dX1rQh6pilw9zrsvlwznT+CEWLRaUetJ0MzcVQKFmj1
M7LGKcWTrlTv3np7F4N2QFnoKzo3DBucM6DFkKqz3U2WsxjGEvAXGXkvT0V+24FSIaAdDbV7q9O9
nyqzZHSZqmhAEDcch/ZjSbTXLMgeb7kf1ORmnzGHVtFJYwW3XJgtnHVxixqbLF21R8OaR79Ou9+7
/A9pXtWkdsatDJRuiiqmDDAfw47pk0hBta33/HmpEWUIDcpKCq4GsnPZxtajpPo/8tDM5mBsoyNf
k0Z0xSHxYoGQZEwZNsYPPytbaOGzf2U2DBy4fh3WLFZ9p9ahje7hA1eagx9T6hXf9/tvXrfkGleY
CruLMo9NP8oPPjLU/zASBfeUXMGWSWA670OZLF3MJExWYxbm+jxJNMzh1eIshTkKP7tO7yN12X33
g8nRNQOgqZyYfEXOxzjS/ybPKaKusXo10EnMpHYClConwjAgz+D4Cz+ydRYLeCStrmOnL1iwtcsG
gfC0riZ1dgY4e5JfltHMZ9nPoZfTOWB9z8D4k4GAIr4hl2cieY3eofYrzI6wH9xslfKwyKmdoNda
DaArk76jsLzB3H1m0vqy6QmUXuQfOnW8JWfRXiYYyVaIKEWpjYbn+uWf6ewJ2hYE0bRL7FytV7OK
SSOVYsPfQoGAtGlWvukAufx7aVLS07NIZEPNNPWdAKWrD6W6TQ0tEFw/roVKouZlYwati2QgKlaG
6w40sij9pEOdDKeYOvS6yU6k7G8JM0PU2EdA0oYjNJWriCPzcuGjeSkjCrNFnQtOUfiZ3VvUXGqZ
Z+JPxC3MYbuA0Eui03yzVNWGxYuIPKiaZ03MoDDbXrqHTj6VDZp0R3vYJXTcqfpzpbIyvXQl+rId
w7JwDcNw21h2Z1NfB6IHy9ru9g/AP97Zs6Thv4z/WJ3AzQAvl4b1bZRjCVrmWkS4/piQ/nS9PxJN
Bpxs9uA7KWbtRJ6DMFL4KkmN3v45JQ7bCBLgPfdGKjLsw8qGJBAW21rrZpHeSwSu5fqxdQztgmG3
pVvnWw9T2zgdagg3d2XtAkNDzdYbW7fW2Mwb1B+uJnqnS9dDyvaqlXXcU62lQ7XpVC99s62b+Km2
EQTl07CvhJy745nE3vcJllzcg3PCFhQMsDnEjpUNQ64Lil1E/M9epMiDwoQVuLewTMwIUKsCdsKz
G2zkrkpjlv3KUCiMQc87EiSzhGUyoZ+gUXAmvthBCr9fDhUABbyy6vBW823C+yUDmVBfghfoROWQ
q5cQfjc1Qu+Cw//mMx0vvJI++oESOq1wbgYc5oxu+yOXOfV2B2pPXOtMzrUgAPe/pQOnPq4I1kxw
hemrSQlq5DnjlMKwG9979y5ZV9kVvRLarKtR7y4vED7vj3eTxidjsRlPumIdYmcYSiQSYtqD3ijk
TMe+Ha/b91OyljnGngskItCW7gdtvdBnvqBBxa8ZyHD/TJgjIRob7ApKdoXG6UUocrfdmitAXSHo
le7LDhFwjNVjuTmsDpBo93gBnSzkYGEhtdSDJVpmKm1W6sunVVFsc2OKBa4EOvahkLqId1UPhvf1
VJDTVr79oXDzXpIqOyZfZ+GZFKQpYBqhrBCzM/1hSzsnN6pNedn/RKnLMI4dvCGBdAMfqC8Y6ovx
lvdj5tmIpncaJJ4009EQ35h93IO1d5dmU/3NKaYI1KyUGjC9xhrafFrmuWGdBL9yIkXuDRCi+AOV
tWR1zpeksrIvlhbKpzrBMi+V5IXfcTqZkJyFL/0Itww6HqQUhtNoeKdRyIhUaHe1puqTgWj38L5k
cOPO8Yt4Za/klArN8HDkDXr9pNmguFr/j67LpAVMJNRvpYPh6qWkqSngaCh+h8hdLXzq+Z2xAGu2
2B7g9vqnxhOeNaa9NKxYKULY1TVWF1OwT3W338VBwKVS7FZA9XUGukCMIvdHZ1NkT68tT5B5HZyK
FPuU6iN2SWksilzcU1o/NJ++93EHOFG4spjInc/AOvZIWVsJcyXjsQaNAfLZDXv+cowCSwrJh7YE
eZ058Ce3EMbREkKVn9oUdJdBRTvlX2vZQ5cp1QN9+tqccTm1vwgZgX9o3ABFdpgIx9U4Y+oNUHUj
DoamEpjNwtSCVLLeef/hq3uxEIuyOPuS9oL9k9WrXO+JeJxsCd78+t/hoPoo1KugiqCAcsvobE7g
oC5YnFZhXWZPL4p5xiaZ+BwbULze163AhHC3a7tCxoir59NwUrUoglbTf5vCC3CNcFIo1nQaaZp/
fEv2JuFn1GKgPAG3snVPnQIJvepMt5M//vpcrcY9SvLoaCKIjmyX11Ll80KnFCNj1L9m6oA6Vgp9
BfFAXuBBu6yYqzaymki3ChULlJ1HZqDX8eg71gf6wEijQHb9HzaGlftMnREFhdGYB82rXM5+P3ZU
t0s3ammgHek9v1uakpzajs/wtPYP8G1m95AxBBbBAIJPa4LSAiMmVpViXh30B6tVsAFsFVy4pkE9
3ROUSnYoTH9Q4uFun+xMhIFdH8ICZCgH6Amk+8maOUNgOGVZXDTEEbeoB/uxpP2dFrl8pOj0Erbv
GEgmdCh4QvWKz6FxnZ5AAD5bC4PUNkqOs7XscHHJGvE60eNL3kglPVOery+ovwlFJqVaK4XtztxU
adlXsPPtZLU2BtGovFq9kkQlACP9LrrfAginWv466T4E+m6FXIuT2OaMJ8AD+hN7VHj5LqwIxNYX
uWUQT4TCgEB1fTVieQWsEhNaMMVSXpWcdNw+2GxGgEAsWtKk/4+ppD/7KEWZ9JmJAI6Xq+rfWkcP
8yw4hadPgpAa4931QXE71uCgoCU5ZL0F3TVUJ4a93a6/caRkAuZhbud2fK/hFmmV+NrM1Tgch5uE
NvKQjtMvuoqmlaXCHFOUVhbj48iY1eV3qVc2zv4pzxF0KBQqpVQMvzk6Kv691DfViTE8/52F5ENB
6pxw9ZBY8+6IQIfvU7Wxn7B66nIbUrVRyMe9l51RKOkbWxv9vQkzcsRfw1AA7Ib4ykbgfhdr+yVP
TJh3Nz4OSj5QDwDIRoNyVr4o+FbzL4ZINxmiG6lOG5jv2BxDCjTb1mlYFV0jFyva29/TcOngwJ2M
9hU/KHXkqR0gf9UdFm8qrQ0la8bt76yEqhm4AwR0cPGozPxB3x+FMNKxpFeuZ2RyCgjoi4LK/IoK
pJrKC2eV1+VOd+d8dUa3r8csy8gRSHKJ1vsxFCaioKWYbp9b3a6O6L9NSIX3ngVBj8bdMfnS7FDz
/7Y4+5fVHwtjlC1htdt+Y8wqzsd4dmOd1jaheLHxkDcsCMmJryiYOFYYv+t++sgGP6zTnBw7sBh/
xvztqWhpwZZ4lRzBVPFuDSg7YNHsmL+3+KdTZC+CbvY9dpKnroBW/SZ/6hJRB+sD/cmX5KXP1bk3
ageHf74EyMQMK0tcWrwPvoGKnAD0o00E14Y4IwG1NFrQZjY0E9YeGvGV3RDfe6YLeEXsr2O+nsar
k2bXOdzbSR33oBT8un01ODtXtkojAdoKPb5atEFdpEmjxy8iAgTVp28xGQ/zxVnkrKqe/6++HFYa
9Vabs3V60Xu30UuM+65vZrHWGCPO995t6EiPk27VWpMSnv/HqmTZ7w0dt9hhDTm7DISx9Rt/ASAn
BojNxLdWNqnJ/LV9D7m4WpoOOYcbmqUFOF5L8oIxSN60PVeNGmqIETFPWy8C1a7YG57q2gXXa/bA
pXLqKxBwb7+VrsTvNV6QQF279gJHyYfeJpcIqMP6zenff77CWj01xP2ZVK4gPR04CcB+iG8YzFLM
GTMrUuejdUGnnLDM+BNoExu1E9Bft/DScf6S4UOc1ZRo6wBIulTIecZxj5uXNYDHZ1ad+EnwCuW/
UX540oEXMUZVpVKwzwhcdUtQ4ShLvbHiaxBD6iVnb3CHXTvrDLrra0ToeL5osQ9jKxmsSisREQtu
+KWKptbfgfuC/SmA2jgVG96/R8xEJI+Qo7C80SGU45maHfZHUnoyLFufkJyyK894PpLe2spUUWl0
hsiOMtX5PSyHBYjfz2gHIxD1SjhvtmlL0A0ipqPAJVAjV9xmoLceq8cguh2cgpFEKraUim0QvRON
VHHKEfdpdPwhHsYUiGn4L2joeGaORCFfTrodkcWtFGqDr40QvJ5T5uZUwOHbrGlx2v/bMJPkmK8W
5vEcw8cN7bTGBrMRReSrioPT77TXBCfwc3kDHOTSOqucAECffndOLy3iq272qzrcsIDlNB+oXLrm
EYj4BhV3Xxh2L50LkzC7H88LHUCeyc3ngcN68PtVRC6ckCKiu0AjtUYSrI1RpcUefafwlB/OEBDO
/HuHqJMvfBo39qDzVpJXiPj5wCwRQoeOh685AUnlyaf/w+dzWTeDA7NU4dBuzXlvAnlDxYeCqN1x
WUa9zmuh5TuvjQsGD7BiK9wlgzoSick0dnG4FOQze64MnGaaqtEhlcJF6qwNe7SJtfaobahypL+o
m0sN+CIHRHK9l9rzRnIrzO78/24bNTwPbc9ueWHjmS7nzqzgL5WTI8mTwNr6SkaabfnuM5fwCKBC
4NfST0uGjeBtBnXSpEQVZqbpkZCNVwOFvPYaZDn3fbTZHJwCBzzWNRYCnUVKZMOjtUCbY76+bxtI
k4ZtE9auCPtTzi2gMmzmaP0xJCu8dR8fQvyjPaMgpeeyMS0/0vqaFXUD1AWqToNI/ySNgXkurzLB
as80EDNqB/jvoIHOGpBlA58CW37cNwRRrtda2ZmvaTPKIINRtW3gXJLSuh3lb4ts42imjASRgaek
qC59dSVlA1qiar7kD+STP3VdKGHA98g1isRyNnoykvxyU0zxGcc1z6hWbwmSiBts1XDN/n8xtgNP
S3pGCyG6vlSIcPysGo+Bs9azOyX1olMy60VCLZ5081gQDtuis42O126WjZaRlO5B1apjSSRStxbx
D+y4dMTPUGi+xdpuvQp/4x+Ci5yseF7TwjlDwfc6XlggURysPu3YHsykIHZCn68TmVGq9wOQZ5tC
JRKFUotTf3O0JQM3uKCBXxP31Sa6po6ERV/gMZgn9X85bYVnrocuxKkzzoi+90608DPPvj4Qm7ny
gkZtTTnUzdkQwPNSPz8wCg5Z5f9Ef6BqKi88oNsq6FFlwPhJ3k9+nOpTl5IBt3VXCT9qN+oinTBy
dHTc8SmZ7el+1rVSWORLmD5yNu37GaxGd0ayFq9TrTGRF1cw0JG/QmhjB6LmBHsk6snScnxTtxdr
h4wq6ehuXkhM3ku0pNa3oWAIQOhU7TGQCwg2s7Jx82UWscOpHYxdC7BPOC8bAF0yzpXS7w9tgcVP
iuN7/b6ObItwbd/dvHdW18EAX9tLhudAs/al79ilxs8nvKGifMwCjNz2/Tuu1q2zzw3kFJ4z1Lik
hIgJm/bX2/zz75WmQQThh3DEfaKZQ+BCb9UzL2YvDgdC0jvh5Hrlf+jkqxAZr3fx+LBymdh/uv2Q
XhchxEb+LYc1ZPhIsw2TAbWpd93PgUBCg7NcVJudSelOyPs4lxjENsybnGLuQ287+jG5+95eKhq0
JOJhdpdIdS6gDTefS8ea2oqM/kNP18g5oXJcIEfPOjOoJJS8CPeI+J3ya5fQiiWtyVb8Bg2gHDes
06nYqUN0VnReXj0g4UwVgZbZvTVPiMcZ6lESO6uTKYbGVgUbm57IxufAKujBPtxy9VhprofKkEir
AV3lvBOSXiSc8TDm5VCGy693ZbafaZepGk7TOjw0CI1Uslq9WO2TAxz75daTfpRgqHy05AlTPgm4
Hrb+hzfwLi3W9qYkUpIKPiiZk9D/EowIoqhavgkhlR+hrZAyUchWIoPRBRPwUOb5SHV6p3iBHmeG
vMrGdBPsahA5BcBwMwnXdDsOVx93oT/pbaEiJJhBZ5lbe4UBHvLm2vSz54XOyl2kfGAyWRrnKUF1
B+J3MCArfNXoVR8Ee/+IMK1C+ZAh0TAgAkLixLsJpBtvu4o5KaYMFHh8llAN2mKTwVSpOm+k3zcM
r8jiXUJL3zS0k9TEfeBtAIsVI9AOi/B6FCN+b0tU6QTKL3vLl7ywpdb6W6wUoiWEwANoKDDWlfGu
cd6FXziOMmTUlcbGuwaWM9OZOIuTmsHfISfD8nMhWiFKI5TdYHdt6NzUpa5APRU9MmllFIdxZMp3
ZILK5rZfNXYXibesO06hhccF9fC1oO3XAzADL2C57zwhIhkWDV8QDokHJ5S9pVjx9j8eNJ4eIOrJ
z2Y4vA4rhGM7cbhLsfl4o3sK/17bm0I8h3PnrPxjz5aqFsMLpMYL1V/8H0Kdg0jTZw/C9FMAk/rS
/UjfeHIkKlKJjhGza3jVGPkDw1i3SLQF8GfdkcFGJTxq71m2Kt/l5EAHjoFv4F1SZ+sEZ14zh8Iy
0RJPgrBk3LpFRacLP8ckBVZ0KZqwdmNOxWEkhXvoRyCUrjC2A3nSL7k4JPkqV0ikJ0mRUAAjhiGY
GBQDlC9KZq9MZpeiwosxcuhbg46a+1S3QqJOGd1k6VxvWBTuLo5xkUD6IhZFmHpgfTJCQ8trY++Q
lbRng1HKUGIIiovmtDnCHQ1WntVjMD2+htD5O/TXkeDITq/meKE7cLn6OpwoBsoFaqbEJ3C0OeM3
E5v2rgtbAzOXE7VcFVquUY2V33f9xV6wuzidOdMpW1b6T6q1wY6+0SUZXvosmoUFIv6eKVrmWTPm
p5A4oY3AV2jvJ3iOZym5UgTM8jUkj3zHJ2ZWr8VMEfNqtVkcm8wQVH/8srIt4QtWhMqLttcRsF9a
fi+mwFJmniUKt3GXm1xNBRffSOfQBowABJlGMjx40VAVQXHdtY+HIc6az+6IIf5j9iRYxO0JZ+9Q
2WqJ1tF9rQ6CXCnZGKyd07te5n7t9dm2Q8/1puoXqqJUJdqEXBASlK5pSo3VM5oHGQd145lXC86B
8kjnuUQhqAghdAPPFS437QfrmJSI5UEJmiMu978Iq1RPP++S1u302uAY4MmVL7mYx7w76Y1Xomuj
/wlYSq/aPohVKj9xPGajwwsooa+FyzaQNIA1QKBH4YV24F1jxrTYWAX8nY+FK7JPfgKDbUDLv9X0
ly/TzkE1fxxlsJ2ZGt+3MfSnsdThRA9orjA24GeXdi/TD+zJupkMrHraGrukeB03/9YZPC5zpA0Y
bqQS6Y623NwcTA2REWuLy2hZ5up/n0LZi29CjE3ooXnkgWyfDkPPLsFV4vlfZBEyb/ptA9vrPo8Y
AIqPf3Ca271BunyKBAE75OzKrQflVoeeUK0MHmLLtIIv7KwTc7ZbGSn77vTs4MYgtThplotCgdbG
mswe/JFeS+lK3ldy0MbiOlfs7ujnm3o9FOku+uEIfG8Qk7cZO7G8YIAP5/lIyBrYsB/w+oILIN11
juENrKdmTA4VM/O5A1kcfYaUjA5b2HF+n/9Va+/c9ZvAwWvunYfVm9+yPK8JLOLFcNiRFukfYc/N
2Afv15IWx9kpmW/QAi/CD7UZRuWVvCibJIHOtK0kFXP4kfUrMBKZC+6l6wTBuByfxThn/UIpg66U
yxmU9BdrPY4aPb8KtQjePn2tZpDLJhKYtH5zHxtq0I9eTb2Lix9SIttOvtRYoCzm28Bi0ZVtCBiT
wjIRy7gURkTmX9nCBbdcftzd2QtwLRec6yPi43vICPFrs8ZOX91WABUMdBZ0cs/+8oOS7ObRmcWU
aZLI/J+JzYTYh3Ds/Wc3VgcSiG2WjpqKPzN9qhzJvpjzimEol/HoxX5xXnqVwP84uZWjdbyV1Clm
f4zh5ZPoHUhMnEcjZZaIswCQEB57/IqnhRf/TqViaply7UVwKi1w4WbLUEV4CDxW6xiNSi0SO9Rr
Q45S2x3vqpKrPYMFe6hFS4/bGSrDSCiMLMCQTUz79x0lMgQ3CkC+JoxRQMXNW75JfE5qJi0Tmyjs
JnzOx1DHDAA2ZSG5xYQvTSsnPSt1OPSMZ8LTqozcFENeIlb3r5SWClm19RDWH9qA1pggja2sohfl
KNg9qN9nHlnJ21qN/t5ehe1COtwllgfHY2ZKSKEjC8jkveNxFiqWKICnxHlK47Nm3coGPL3auxlL
biwxBnis+YTkA9J88ji3LcGt0Ws9Wd+p4YPeP0AyR8Y8qMqd5SusgGbANgAiErVX6V6EQn1rXNCN
FkqRbit4nX5JqxzFSd5qMBf0BVw7+hsm6nAi2n96D8azVRWNC7FioD/dZUX8cW/VmIuWcy+2Zzm6
XFNTb98pvWxDWkp3f3Cd4T1DFV/co+yZFbGYUqtuZOWABI6NoQX5VEST6dyfIBDRF89oWgH2bAWt
6WYHkA/XWHGVhFXR+Cytcl9AZj6gY1bqTDOH7p+8rLegLDTAJLIFstx+oPDvqCwVlrpr4ZOIgmzk
+YLlFgjetugmPGGvCfOOkCH9/+IkVkXEobRIZN2jk5JqJDTXsr4rNrNbg2kLbwJ+sF8PoYtwWqqU
fyPdwJZpyrTAb5xsxHlhblXpXt9t9LTDiDNKA0RR1JH/Y6LafrM4Dtw8waDAd3TuaAw2Wes/WT5x
FCp7KAfNsW2tvqGtMO0TdCyUifucOgy8uVj494wF5Z7C1oiJEcFJNg7yklXRM2Oz2i/nTQrAFwtf
iXWIYK73tJUZ2sGzzidjSFH4lELdKmEl23HfnWWEC4x1004mjxjOn1YAMb1i9zb9b7JFu5Sd+yST
u7PXgj/UACNYaQ8cOr1YaQ+ECEGEaSqoaTEbgDh7o6Hg0OtTyd6H5xPIAgrsjqEJs/I579MfDCRh
le/q5Us4P5l/7zhkFFgY+iHWP7u+HhZatzGBrdAHi0aLBQPMs0hLuJwg7weNCr3SRPXAQmjxUyHs
czZh5BQFiI+xbntKXpeWpzmEFZ20Bl5pcsUVTH7m/PZW/uLE4xmdS5qWSUT4c4Gd58ORhxD3cFS+
cTbyhUaBYlDDC4GxP2gbug9NFSHesFFbt/F/TPVfOFv9mWfzcqukYdVVPdVZtQh5PMi7XK8ne+/B
jqJcMKDoZ0bVH4QMYhX5JQ9h8tBHg3MDC3tQHFKQ3t5DtKNsuiJ+zbj7/FIQ69O9oP1SqAL1dXi0
gRHXFODDbvtiu5IjxWJgZa6/ALNrxj1NKGejWXf8Z909M3WjkPBfaPqzeYvKK0M4lXSGb3+6CFIz
BwVuJoxQrHQFHBvKSmLzibBz4DSduLEINXiHV9+Y90fyBplfJoIKhUKyHujuavhGllCarAQLelG8
WMPw74VE3PL7r+73f4x1yGnF7HITyeDGGEcrJKp1gxcHxr3YjMwNY+aF+dwyfRF2pT34JsXMmlvn
zLPtT19bSZl8so5zQhsatsYjpGXvWB5/cJmdKkcWJ6wUDIPfT00TE2jXx+Iau9jJpndG7/QTwRnL
7w8bz/V5Kj9YmNFmq/5lA7mUQtaZqXr2NlZH7tWULUyvjFSEo5k6JbXnzBqygNdCZUnAHicGyTw5
knBNYui7XACChnDuIcRIzPuXx5NphUnE68IvIQpqGzOZwAd8jkf6tM4JvMa5ynJ+vVRXby7/ZlSz
Q+MKxSkYRf+3Gqy1UELw3u5Xjb1eXog4/PhWDlcxcc917vIL5hGKXwsMYdFC0mflK74L7ukYfnN8
fPwG+J1CXOJSQeYobf7o2k8Sjjn9k7h1uYIXyuZs3qr8nIeV7j+TLFnbIXxjsijW3bQpZ4beORP5
rxFZJarJ/GWaBZs44OmM6Ns3q2eLI3yDAmnT5GNaX5ictqIbse+oCrgODpAgirj3kcvEmJGUNvJd
o/Cyo3PDM3K/LhJlBt/e9juNF0VCzob6hDtTayai5KU5DVJMAKRZ9x8YF+ih0lXPGDv45dJr1CLx
SaLy3EO4zHJVyPF+PfuCce5B7Xyhvpu9U8S/K5K6WYdimMLddb0qCk8BvM2SMt+uxFYvD4ReRyft
7wcXvwFNq+IdLzxLGz/FLjvk25ENYjonWVDPf+6bEwyz2XRIllfn9pEQjQ1q/m706RGGqhNCtNVm
W+3RoxydBT/NvPaBpN1+t7Zc25pLTCh/frkPIqKnZC/sqStJZAv00XLfnTmeG2+m4Cn1t9ocf8vT
Xr9G0N4p7HrXSASD1dtvD/ODDvKSxbPuicPJrn4hpNyaKfN7Bb8L8IEd4mMCpP7Nlmn849ESX49x
OGcMflfjF9szUvZuFA/hBX7zii5XS7Oaugq4QyTwF66w0m4QNifzdDUgrashqfej6PXy4+fUpye/
H1lCq08f2akd/4E1l+/+fRJ87QEX4tCJVM5fsue8OYCjK9zNJpIy6l7ZIaYR/ZEtufs9yUXcB//U
mwlltzPABpIaquJrZIFqDVxzgkLvtaLmWasL/XyySI4tUJApgL1l5EV29snKRiV3Xc3p3AE3B36U
jbfxFG+toiCOcG37bwppfq1bqWXFAc3vupU2nu/IzgHRq5lX1wTTLReTfV4Ub2va5w3LNqstQHEP
zn5wEMZOeyQxEPbEVluRrM1MAOq22SE+ci7DLLLhuLy1cZMSyTf3Q0szH/aL36UYZCy0ola1L3f1
F9DwNHiTxgA8Ui3Xt76Ou+KWMfxn2PQE7UJzB6fJxZGFVS4pnKD6zk33qrFJ54Rjrk01wpJQvQ94
9IvYpaJIAGQeNitEiq7WBLMmUIM1vX2MkPcGanFADXfvdbKnQZgnOFhUN/GLUjZyXsRWeOdUto9v
NcWPEJcupHMn0mUHIJ7bs/UmVO0f1EmRYQBo6f08Fv8WQuSe/R5FB58xX9rzFBAdU7108c18/ydY
8wzb/cvciLPJwi8H2FRgoEc1/rS6wpb8LommusuJnqw8aZqknzQo1eb5n6Qc+D/nbdZBWtn6A2Ns
VIxPopefPcz+2/cLi4S7OOPNUPiNmxWz+KlviIJramuxdNzN+ps5euLohF1YN6vYvCC2OxJSl7JX
6dQOW6Ved1HCGthIMlOyiYFFTg8+kybBUw+Hh0rMrqOSTh2AoEZMo/a2PjFJJr0IB96XEwgeVp4N
aMP7kv7G7C4gMakrh/BDMiFWj+lzJRA5GtLIp/3iEqpxL1DtklhzAkEdVxunaOHHoCKvAA9EW0UX
PcMXd587oJ2AYzJ4fkHnGKHedzS4C3n26XknOc47RP6LqOgGQdOE2v3WqgEKTIJU1iTngBuRkg/Z
Yk+kWIGRyTnivE5k2KuBTq/YphBxU+Uk3kEjfKUmRMVf/B7O/jZ3z6VHnKVd8i3pirJsedhR+v2v
0HONnCC6GKBjOhyHsO/e3ngc5sBHtCSuKoNVtgSCeJ0jPTx1Zryvo4sIozN4MIEeZs8jXAy5VfmP
mKVoS51Cu+Vwu+GKlYHqv2DcEasuGaP+6GyOYWWmNpDq9MIxPPmc9ysaM55vRUzJIcYCzoWNczzy
5j84MXiAmOoOKBZane81qKqPHIz5LOuPg0OmBj5Q7mG2E2pIRyLzyDBZfC/vP5LRPY7Fir771cmM
fznRMhfqHtLe4Tiu8ENtG3kZO+zAyIOqr0z3Dnr1I/OZ8CkWoJXkhy/jIReb9rhcUJoo5NEHXTk6
wr1rA2yX8g5ULd/0ZySixahVICRngreJjcZNKsShDQEESeM6LQ1PxCj8sqFrbX7RMgHIcGb9M7ZO
xyHIzU0Nno6NP1ih8opRftaj7xnBClRYCQaQ5AMXqST7JFfClcPZ7V49vKCJhe2u7VRX3Nl2J+e4
33eMLnWEHtuTkjkVze213medqtffcG7ATsh997xUMwuJeW6AsM7Zg1YFUodNkTG/imSl6hNb3sPu
vyBbXH1Qd7fqHWLXA1pPks6sqEmUP3WCXenRhaMa6U2lEYsShsrM9IPf3CAI8L+RYlatWq+FSKZ1
rUTZxvlREZaOHSIjOFJxhHMilFmV7h4XWEz53KGNqpOnWoCax47O7lWGVnL7ngjVCzqiy4D1gRNr
+gz5kFb63QE90Mr7uEUsHBi11IXtdt+dJvWkXJQjo4tCCEnCv+0wj5II0zfgBkMu7IYV7Nk0oOmg
homlkR/houvEgiysMXE/u1uoeIopj04pQwTpVS3k9/VFjnKiw0nLitxUSrnbc7u57lXZZTTcphqo
e3L5tbsNgr0b2mWuufm+h22Mi+k4BbsCmZYX5DFx0VMz+9ukyTws8eNGUlkHKB5weAMzpS1nJqIP
Fr5iYVRUYctoBPzSpQACwRVZoRItwP3B4zp2OgiIxLNY2QxG8MPgMruifZI6UFzQ3O8qSKzpJUbx
wC7xxSb+w9yeYeOOn6PVQ0PS+fqhmzJZuYAz60lzZpjzBXKCfpnvRe8cIXruimuscG62wnkgTWNw
GwLT67IegRYv+S/yQS7wGlCvkDr1NbDY5ot4vpsBIwcl/g3Q4auCNDu8DuyS8l5TToZhNveEf2TO
xCC1tjqHg/PxNjll14rgYTnXC3QQA26dCLOYJ3GUoLQ9Fx0UeZrFBaVhLBLApDMBOE27EeITqWP+
W2ZCczBcuEqT6RoD1H14pMn3rXo9iXuPmKKH6snwE8rPU4sYEIBECaI0haki7kU4G64OIeowq+Rf
64/FXRJT2ClocnlqcRFWidxGWn6HBDVYdBxBwvynVmHMy+iUS2/iAKeuDYy+1VbTwhNiPak6+Uun
do3qxb9Fwba6E2Ru3Kvycru88e7xlc99WYtUFO38JWvfe7dXq/fEhRTy95tQbaQcd3jM8TX/ZMxF
lx6VWbbDsG8BOLSoaduo/4KWsNdQ7oeP5jlxU9DpCrSfBI5YuVdy1ohKx99wSOdCBW2XMuIe6wIH
G4W6ncLUG8tMiw14EqP9AcFny2PC2xUzV5ImStM0lIA+ye9OsdW3skwabGLevW1a0YF3dL+5pxeS
smPnUFPe6+Ng77KR8HRSegD8LM4AzqAltwrq2FjqpCiLZtmAdXbLsWT+hTnNyLNDQzPgMyQ3kRhH
vLWjLNIull+L7WTzMwO2gn+v5R/y6FMOXeUd+ZFYDb9VZ79CX37B5W6HcoQSw7dTccrif8+77r7J
qTPjpQPS4eCplB99/wAARV8aYcLrFMPYb67Kb5ugYVGvkN5ncbdABFHneHvmU0sgrPcuaEhyADHt
u71nDFiSiLF48AlJ1lvYF+ZyqEDBwFklJoO2medPO9T8kIGCJs7ckS8Oy0H3EONJyfLbdCAN9zyx
9CcU+1v3P83AV9gfyTqDc2nvOauyLGfY1sMxtzZety4/9RpCNxM89DehBea9vkvjONbGvPt0hPEw
g/LhV0KIXkJs3lGlTYsaj+bijEdsRWREWhggxAxyfkbnyI+Adn0pmfoVDJHIqROhGnqBslgelMv6
yHMJlEsrn9etVpUEoToVLQTzL1yW13caYwxshQ9D9U12q62IG6DfTqaD9VNE7c+1RfFzzZXwD6R7
JyuurqeP+MCReYFHGZCYI9tGbDuyV73BB3oyLtcF1y3BWMWbtA3jX/aQzAXoYOnCTzjGMmv9tNEB
LhLmIMwBX0sheqD8xbWhWiOeTR6dCfbsSRClR6+K/1xUuX5JT5l5SRx4CkHmwyftoG72KpzmRCC3
nf/AavAK7y/f7P9f4KsAoLxUXO8jI/8kG1li94V94Yh11qgJJJQGg/OWTL/805/yN+085pnkOBpu
dhiVf6+1L9GUMm2bMiuJYnSVkUI5J9xj+km+j6WNdB7OyNmQ7qqOwRUXO6dx4fCcZRsu/npSH4Jr
7N2ff8HvzY01aEa0fKKOhcaBfxoPAaZ9IY5YI76OKzQA/s6S34c0F+zmaWLT1pQVL1Lj2cFrsluQ
5dzXeXpe9KyYqm+4jxEHp9a7NFsKMScLiU6spaMbnZwMUXSZHz2k8QHfwDE/cmLUcZQXiCroqmh0
sDt0MH89NEr17byLAfb61h0gCJEjfxkrsI9EJ6LCp6XrCJE5cB4g2MM43GzOlowS35+uVX+e+3RZ
dg1OeYH8k4XkUZTXvhDbpULpzJ3OBYbjCHfeuWigiE7Lryq2BCN5NR3Q6ZAwkhhFqFLS+FnFe9iI
MslYBEi1X5gjouEmtiN2aNxRlMRCAguWC53R1/TtUtP+o5P3khgk/DCU3RTQPzlRueUc0LzfDEtA
lzgDhe736lsruxBehH1vKEjv68ge9DySHBlr2JRyC38VGxaBTvPBTINl5PeonIwMTd/VJGdHxXvI
6Xnjj5q7/4lgB/Aet0KKpPzMQ//JLCwIGFTBC1ET/+oTibAtj7Dm+GIZzVS2FJqMeHxEPuiMNRTj
BdpwIo3xwuBU4+C+43d+DyOLHhmJzlWE4QpapA8hpRZs/TODk4d3nBysm0rFEvfIcIg0ZA6ORC8T
OH/D324rB84nP2UCov3LtiJQ0N29Wt2qIykVooPGVMGDguSZSsREOpPWfsrVGD520NVPz/kb8rXn
56ot3D1YyRHmvWD3Sry//+wJFFAEDATkASNOHDfGzSq4Wc8/8KC32W53D+j+yKWkOks6KH2R66su
mXWnIgJciHQeTPiZStaaKmAlrTS3foNKGPsprCVSNrLVU315W5aLzGuynPVTXs1pLOon1xYUp8pG
DN/aq8i1mCHuVFWcjzwQRPZQY78jUIgBTPXaY/ZOYDrfbrMAnD9NcU/7Sq/XfzbXLNhLpFVVqJ+R
zjjco/EpWsi9Kqir+wL5CZy0dtqcrCtg8iLVF0E/s6WWcBojaINZbp3E1huDLBAU4pd+FRgVX/qy
nLNlOKqUxLs5zrj3Uq7oJzRFuqhAUZ+foeUTQXJGEG9pE+YTlyf2CguuvndtU12zaEz0ziJTrvje
uLqUAdot6QTPFzLUGXmx642eYxK21pBbsnB35MV7c0KqCGbhcp5WYHhqI2enicBref09YJI8cgpJ
wSGdRTsvlxpYT3CMlLiS4EiIhKPRZRbevWKrUH1cqsYAQwsSXwPNxVtFhDg51yZjrtFZnLYCASH0
wpszLOJYQEoSovcJS0KHMbQoe6atuze6U47LrqXf0N6Y3aLTHQyi/TmYN4gAAT7rDpR4SV7NJgim
ZoZ0ilLvfVC92UKNzbC0UVY7OCXOKlkkGNjmc+hSLGzAsklddfxSMPNJ7knfVozIhp74VoQO39R7
gAdfXYTmw8ypIkaZZBPX9kHplJs3+la0c7Q+hVPu7abhyLilxoUfdxyMPoUwe+nwnZ6KzcJ50Pu4
g97ypykX/k8gZOPnNRkC1TG6abj0TPF8WlVCDKcjsHWI0FjmFGvXbiYZDq0lsJRHWVuH4f5bG4F2
T9QPPNiOdsRtfYwrYRk3yVy20FgvWr42sJmcS9Pz6r6oalXVa3VUWiztHSEN6v5XulXqNOkeNY9I
WRw+CpZbaL2BuY5xYYZBkd6Vn2X3ip5vFiylZd/+YwmeklOY/Pkg62xQDZKADS4dvKlLViorUsw/
tnJZKo+V8YDVX2jrwNqJ8vGF8GThL1W3WLMGXGLFEbKdlDi8Vk9SKafx5ZD7Hi6fqOK/ntzSsAW/
Undh3xibA5rNtYqfxIWYfLU/6WvC58WX8vc6bOJI0TLGOynHZM8pYnn4hESJO1uFBgdxvXncIiW1
8NQRT96mxNarXsM8cA+EQ+9GMtN5sSgh4DwKn656bcGWG+ztXqs+s7YuFj22ofGZ9XKP26+p8EBI
SN4xPkfLVko3jpsGxeaZxnSJyFfRgxNC18LWyKBtNE0YxFNoq6E+iHX0lnFsADzWHcM+G1RYx9EG
A9bFHCBmRwVkLg65xde3YsYRiyDvslCmIb9krD0H4cTbkKGxbqV4/UUOgKfs0xhXbNq2ic6dqETF
NPKgE0g8lyPAio1YmWYridL+J7uHrPBS/fwkdqhYfY2mi537Cv1kHYRztvDxF7JWi6+PBqV4bxU3
p89UfmBsDtXk5RY4cpeMbKMOAIMhSQlFf6K7DiUEV+W3Cz7j1OfOTGlw0xmEtN61vYll64RYP2IZ
H28OspphMMRoGSGTm+JeOvFsVSp+grbmz4NwLspsUuqgPgks75wcb7tFGWQRLFyzuwiV881tuI1N
ta3IQ0ZEzastr7CglGjCuQptv//h8yqw2z3H0QhjXDgXBR21p4T1SVaU/RfPpAM7c1+JqL5jQWj7
f54qIN0z9tPJz4YJD5h/qBEDFxchPeUyl9h2hf4e67gLuD1NqMSAdfSkg+SveGKRtM9todqDOxPL
spEMVfUt+e64/uM1LhyYMVCvn6Z5/fxxmgfyQ7FuJ4wyJ3CbyJVpMy+p4SMbXipNR+ZnCT4Vun4B
X5wAKyfFN6pQ7CjPQW/5WW8x6fNi96cqmX1ELC2s/zhcbqqWCyDyw2MBruCGzvpeaYgYvhOHxnuJ
ZUrF6+KtyNAtbRt47PC8b3bfPEEppZg/C2akMWyMabuas0QL9ggvFWMSmgWaxcNGzsM65Bhs6Pns
e9kGP6K0DNuD+WI20pfamMiJjy6viDtaciysT4cUdwwtVXuiOak7O69WPDs8g/0lWKIBYpPVCWVk
8eRsOUd1kYrS9SEtqPps7uTiE6GtkspDx2QOHbIJE+KDCKNQcGs1Qlp1VfLgdQwx6APexh4L11yy
aov22kCd8PiurtSS1+ScFZ8vHdzCXqZzNURbBFMp2+4wlNoo6Cd5+idlQRnc3fpQq07TxFdATwlz
UEszZO+swRzXghlc3nRVEhZy0fFNtWws6LiULRjJ6xwOWGCFLlv0dqzUWaBl/4VxU9+3ZS6yeYTh
halOKX4sVTGsx1u868BwuNow4mjy/fjkNzZvwMT5OPqIvDRzFgyifR/EEq2T6u+Gpb9WaN+F7Yio
2StRk4DR5utOCy9W9S0+P8DaSVIn8sl6ug5IS7IIdwW3QTSncDJ0bSj8tYGWJP15yrN5S9EzvYDE
kYAw+/2vOUfA80Lljldf0lTjT6qrCBNizzVyQ11RhMtjnUhptR2HtcUckgV2hCEomvPSdRQaid06
ru+XRaRpNVuo2a5yTY2Ek834lULKG3AFEodGpmVOVRlSsf5leW2wlJCtiK6TryOHZs8vI1mPIwMl
Gc2fLpWifDpU4PYf0t1NCmJwPlYaHU+pMnqEN0ZCCazF4xR/SdIIr4snWJmlZl2x/AzGV0mGSFDi
ge6CPJuvkpKQbbIvJ3lvfybtLYhYpPpHUd1J4db/aVEmV+m+6PlQOlCFy71c6fSw48OCbCltIj9q
Pz50nVUO/FJXiHeGId2puIWCzbETmVN+cPA88k09WPBSFTUJC2vCq7bXwe/SnyrkqtDIqzrQUAxN
XUM1pfqMdojh6ElTTAmwimWstzWNZWUsSy3ISu0gIACb6LJwKQBUt+vRo7SDD/Mw0OjkgHNegzrl
e61bxoAL85Ud2XlZdceMwJbEpa+AVNWiCy8rf5dB4+t4A52AC0LkfEZSqc4SP5Tgb7PWV6Mz672O
ZYrS7oFoJEvmMVdsllfKGILO6lfR5jY+TTNOAu5X/53qY6YVv3+9Q3F1d4FBiadaXwTjCmXxiddI
4wCQlVmjSavryzOXNKNkUAcBiANtNpeo5EUxqN1MKn5eO9aOG/UsyXXavDWuSBiIsMyTaIv8MNS3
Oqwk7aa7kujlWiIRSZ3N6gT8IUBneJqv1qX1rzg88EN8PmPaVWneZisiFgcRJy/piBfOeqAk/9p+
01XhPK+owVExoCGq63W6FNN38u/ox4e9wMCmk1jhWnVi7nVHHfoEiUAuQ2EjoFN6eAeK5RgWg9Mz
hOwuId/cZWS2x2fHWY5qcBpScOquFxDr7/2CZw46CxuqYmHuBdYB74KO4Tlc/EGcmze1geIW7car
tR3F9rR6df9x0cSp43IHIpY458Sts89gNKz7SnNp4QrcmX1BaMZT/rOeQD2QansRrZoZIb73fH4/
5ZhJa8wrRtNbCaHd+4bPEEMz5VlO1S7Q7xCcy3B1TMFGeE8vy55rmWWZlMeC+bplxW27dW7M5ujg
JJUQxuOnMmUNCIfesmS7FGZc9jNBSJOOLLQLku7mXs33fUQhiP0J/tss2h6Ia6hXIxxe7qa2tgah
ekuUwQEAn/oXF9CBUxYFD/Dw2Bak6nU4nCoWaq7ZidXW/xY50In8MAG0fkxg1WBSIhdwbVkqQWxq
xApBydy7YiiiS3kQ9RryzTk8eAWwY0T8eEOSxjT6MG4+sDUURb3BeoGo8IAr5kiNNXCgI1YHWFJl
WMLH2mxJyO5sDt+2zGYyBikh2w9bB9I7yo8BTLOluUP6m3+EPmySdUWS8qpWOaI9Tt7jdaEvVh8s
ym9f0cq9G7WvGyEJDNYSZuWbb3tTV8IxVvx60JS9NZnb/yZW0+LRwaiRb/032r7y3fehC++V7kMX
bOBgZCiBjuZCbo9lpj1BS0ro0qkHwK4+MmSpjAlSSeHRBbZu+85N7ZPr35sKW/I+ErkdhXU/gV0O
SITiN8FvIv2ewPcXGA/mvK3TpyUnTKVGAu2547rHO6a6VKHIGR3g2vlK/E2cNV7mPUeLNKdmEH8o
BJCpDvRsjfnYacNHWTgXTchHftM8KkvijXZFuSlmdeQi0o3Wy10u7NA8h9oIgtgPmFcIY4c/174l
BPsTdRSj4AEfzs5TdKkjNBOC3S4T3NAWRmzzKGbd8x5LhG/ViPjGxMYnYYz+H0rGQr8sNt9QAACj
kocwO7Wv/elGeZEfaPTKWGRDrpsal0/oPThafyp9n5PJASlgIhziQHh3lFWorYmKb8C03AtCZ1kB
5P6m+h7ku6RxC55XV4wmhRjSvzrV2HGuzoQOc+G/5yqwcmoVixLR+r417rZWWbKUuv7OdQtnTC16
5CqN1SE/x89mRFV8LTVyHVq5c3mQf31QEd4rq56aj2bIn1G9TDMr398/qPwgXLFZ0BjNrrbULfbt
Vjz8ee6v4uqt8FIEzcWSUsYaUWPLy3KxI5iOOjRr1euxhTe2BZZ7olyb9Sq1BEUD5TeL6uEczkA4
ojA1hfNhP1lVkdO/XHCcgOL6gm7uJKKSXf0TYsroquNi0V5u9r8ZS4KmpYfOr5pOsqnh+V4IpyhZ
pRJm43rcxjdjW/SRgVyYtxVwLz3X5xXtELU6ZJthN0rRw2XIqGv4Ww6J7fKCK5xi38/8mETZbKN7
RMyocWd08Id6m8iFo/t/w5eJGgDz7+1JPET+Hm1+Ce6hRfkEKMA/dCoDAEzyqOAvkSlyM3bAo6vf
FMq1QTiaAPXZefEzc4HM80xMfOFRaC+kILYimF1Qn8yQc7XxdIlceN42zjhXrlgHdbp9l+vuuddZ
STiTge+8hZOFUnQID0LvaW1EfHcSxrAlq0n+7L6uUqwaDb6z/BAoJhCAb5PHRcMCjoNAyztkWYDY
lec7dOIfJp0vu4qYJsBfhVtcABFOiQVGpZEaCEkPdWDH/vDWes0u1JX6t/rKJQ3jXmxuda/cRbnX
Y7H8oVcRupiVWrDsDJ3Cr332u5asw2/CQBVhkvT5hENcfRjr1kMNYOtWBuzUp+leJeGuxtBDzZ8e
aUBi0K7NRLO7R61kKqAnee9yUz1KTSCqNCeyNL5U0V8vovrA1uBnK1WvkLdfIUtn0QXWDYaaU2zs
Oy+3AjVNgQSDH4iptEv6uGwDZnBQ5PI5Ag3lDv9xmUvPFGTsxmmZa4MieH067itngrscO49Q0UMP
wwIx/m3vZ3PytoHIRpmb9F5EDj42sgJrrOAXXg6qL+IiWKcyx1KCYHYeEjl3pP4Y0/eyP3C949YK
Gs/XO632miMYQ7cO8mgpcsY5DJcUiEJykgE2L/YIZTnWDII7Jh6QV72dWzaN4/zjJeW6ADb18Jhl
ZPx+timgSed69TEZ9haiDhhR8tXE46WCZhEKx4Tgiaxp3KTe0diKLiuDMMStWpkeP5oKDBPXL7z9
ZFpA4Z5FH2RF2m9LZwQ+0RB888yA3mxRIkBqkpR6mV1Pb3RT0ljBkgU94kskusHn2a1GsoGtfGef
aHr4z5rcvayE2L+gIQg4YKjOPsX9TSQ22TpDv4qOPX+Ci71RLFqto+aQLuOn7EBeL37zBonqVsRs
1M5yt6VFvknhqohdY8KUR70fz1drFXV8+3VBS3CF3zg9WA+Tx27k88b6dQZbBfNO6ffTvEL/052N
MvIhCs4CUJGV6onums+rQubfyoDlhO6jKJyBTBZqI64A40Nb9UkDK2Ttc8kjVCVb4vY3hDt1WTtv
afTihH5ezkgw80Y/376KsNrAiAETFkOB2gJaSEMgPpcPU3LAxMRYNq5PEmUkj6oEtYCoCTH41jq3
vZag4ub5qxF2bTmkIsANCGTod0EyAOpuBvr30ckkdqag/m+yBGU+TJrwODkpUTAT74UScW76PTlv
CETjDGUtf+kgX/FhBWfXAroeIOdNbvl0q0LN5D+LhOC312ObCrBA2xThjN8C3q/m9tSASNX2ciAJ
cu9n+9mMT170UB/ixiPQSmFKEgXirT4+SN/bymCbS9oetlmmCSLjfkfAC471kC3lIrz82t1Wk6+J
k44Aha0fT3f64/xLqh9TcQ7BI1uSKbyMNhKC24aTvxHZ/B9OTXgS5xcCk9ZrSJXqE/i3G1DyM6hZ
mLSu0GaYiVArzsztlyGtyIJih97GSbJormA4szOMh9m8SxeAOR5u/KBgBo+rODlV7m3bCyQK/c7R
XMMClM8gs9vghMJGr26MzsDIBVvIHvw+kTsSaH2TAENHenD/dQ9uLiUcUFuyxcmg8Q7GT0GZj/Q1
IzAxKBpCE70tz1ZS18UpMOOMDHvHk2mmH7Pf/JCcTJI4mzCa+mPIbE3/ogKafsfjcXcqhb8L/ySJ
2FWonV9VHOvvrn9mwqkYUvssAy2mn5OPLOHI2HtDob5n7Zttylce3UudNpypiTKOwArG6wbLDTDc
+jKXBHZ3moDeldwwJdU1H5WavC4RlZwWGx/WA0AF8ScfgdcTzOVo6vTyAam0t20SICl7JKuJR3jQ
8Rhiz88x11AHWfGQ5eOgX29trz/tdC3z3cnNs+1ayJAjx6AZS19BpAvgWMDJ12s6hNwGUe2TFvZ5
1Mq0U2UAmI6iiNCeMGackIB8Y7UCKD6X6laWg1YXdZANdDpPjirgWMGlbL0mXl7DpwByYui20IZd
321XR0BsXPLFH0GpDlc0J4m16fsCnt/t3d+BVFWTQUduOWCU5qH+uZfJVbQESud3RQ99MmhSJrST
1E/owS/7WhUKPwa7icOdPwa4EaxhGF1lSHzSN8W8EU0za56MMH43AH0DmfUUQmxMosXigFznFohn
zjQGZNcwKYydkx3O3DUWQkMTL67JjVHiJpp18gHMmGrR6B6PhVwQbuAEQ5/qCMZpyUBaYfkGsrzY
Ac1NV2T099jkLknQVr4y/AaJtdmtpiz7z3myYUXXrinlU1gcSh5R+A8RS2Oj4enr4DUtHXY0GGQ9
oppDs8VOP1fIPzesLzXiyAtNCGcRlOgkFMWsaU+ilRuLihJnH1TlJ68sGIi6MYj3HS8CEMvukE9i
dRdD+XG0LslM/7DRqUY2Wz/Fng6zXINgR3AnBrFIDmFOHQMrIT9nTfmDHRIqEMwR0RKSnogAfGty
yxxknVseHYz9FOmCwVpPg/XxErRCH3rHlVX9AbQWt7yZRCO2rUeTsv+0I6Z0cjLOd0mLqI2LjGRI
fGbUL/AjDYuVkk5yxn8UHSCK775yA3xQAX102yE8XGBhsCSN0EQyVVwwsa3wLhTz+S0NPsXRmDXp
qweiCArWlOBiX7ln1vOFDuqnEFl+B3RSDgwkb7SSuiL+QyOHr96w9Tzu4FQ7gMGiDluCF9twF6Cs
+URpWWJ1TsZimBOz7YspccP1nQeG1hzP3Zpf/P6TvYJkkR9cesHo94AH0td2gAat9xNafRZTcIOk
cutUMtc5hbYaymDOpSy8XTaRE19Yu/0Lkb8VGX9RuLtO0W1/kjWq69mjROaabgCoS8XCz+iLBcyP
QPorLIjdYjE91RT2MNtKL16RUna/+gk1NH843b3/vqdkc1rPIifSgKmpWdN2XbBQ+3XdgVZyI3jn
VqiMHrAO+v+ZuwvcXX6X4XlWG+yX8Tk1Kzui0kOeUrttGKEcQC6GI9MRqG2tLM5DRrZZPFpY+n94
N20KS+2u4ZpITLhU0bf0lct0zVl5SXitosHCb0LR+LIsIHt47NiFtPO4S6PArKnZUI62ereccrSX
AdWiyZHa74nV1Pk55NfEbn809/vZM3Lzuqkc+T/LeWtHnKqv5rud3Ir4jIbC0H/pOVsRekuZNfDU
o/6odO3yb3wLWrS8eQsKgjKgW0IR/taO2TjOQ6j+Ctw/J1+KFFTiqYOy36/SAWx2J7DQgzJJfkoa
yJ/8D9Z7E/GCxqBBaOLWFworfUViQSOEZm3MZlj9+Sz71d/JrY+VixavAqC9dlQu7tpRyPHWaZox
aQkaZsrztiMFOJOUKj/OT12Xm/d+8EY2E2pTKjKX1Yi7OJu9vy3UCHaG23iOiW6zg3WIVFrpw3fc
xa7Jlvjf75lxLiiWR5kC50Z/j6LJTlMjWU9oiWkrcOXdz5j/bupIr7ftQWq6NacN3JozQRhFAG5x
kpfm+th1sZ0JnShPo9k2nTpzLmqm/LBqB+5J4168Z3Eow+xsTqZ644QPkNExOASro2/24a2SXpYQ
wy1Fv8sttG0clGCBufQ/tvdLumj6k3VtG4z4fJ6wwa9xkjZT8mvNmMcsnry9HLMsI4DK34aZJdg7
N1eZHvx1qcqw1e9WWQ8PpOoGE34IJhHds5fC6Tfjayn56k/plRAezfH4l0AkFLDCB1b2KpiIk8pr
bXF4F5l6HCYs3TdawkGUPeUf2VpHbcqzdwM0M+Rmivr2maHVgda+lj7qTAWjZvd0HTKHNFC6wLxi
xS1EDWEsElBARcaKoPJ3covKGdczhSZEDL2TRjuUyenQ+p4p5jIVrFm/wPkEY6fQiVJw5PWtMPU1
dRr8u3eR15x+vJdH4qazsybgh24Bl4tOfvSLeYLF7Auc09J3u4gcsVEHLgMNo/OdSar7nTTIMQC+
orQfzfWiTVAXZqtnbvg/NQm8lV4qJal9LicUzBOfxCXaPP55b58Ozm0KVWRk19P1GpicTtBQCBpr
LR2Bayile0wZO3bONISMsuSIo4n2kdNhh0CedBN4xvsCcbDp+kx/tyfg0bsTq7fLIF2kYXWMEdff
temuU/TvVoEPzfkf0Xt9DD49kF5LsjCaS/zDZFoYMjq1oOCqRIkpJPZLNN+qy0nKyvdQzJcD2xOQ
bONSOTAut8lstBaN+8Z+I5Zm7he51owp26D4zjsxd0ZdrEGYLkzUAW/lTpcBGYQtfAjeMMBBhHpW
AdX+dn8osn4gNA23jaz8VqEtJaH07vquCujtTpOknrQs+2VPfsvd7Dglc4bE1k1WK1iXBsL7vPYc
ylHMG3rqwecp7CiAaawrpW2wxLexA7kh8+9i5Z/LbWFGMDepDsIQZq3BoFYfE/Cu+7DdGy4J9eRc
k2AW4wBQHm7XLZvWQQSxbgnAGuRKxEhy5cpQvgyRjDpVVpEqW5zHRT6cojThLAF/11xSHwkY/ANc
135l11Tez9e1c+/QjVvq1VY1GUmkYn+l0rbKI57hWWniIQl0O3XGnDrJ+KonOqB5U3QEjqD8SS+X
LNMoIBQIxRMcm1tCuzLA276PQmzZV9KK2Zh7HycEAj+SU104VzDAoqF4RC5P3fTiDcT2Wl4BbHjD
kCGNnC30/GzcBdqgJmqmtf/J55NyjHa8VXajAAR02rfIFEkIUF4tWOA2lo9iC8SPVCRjclX84niC
coDluQhzCa+orY+81wfLKWhUPWFwB5zIiPYI8WEb2C+n6GoBudiMy2PxHv5UOuV8Wulc58irvGFT
oGLqa55lqBQGInAWMF3DP8YU2BMEvVnp9JDKFn4BAo683zCjK7llT06X3AxyYWcNt7GM78CvvJGR
yoVO6Dw0pKBhf5s8XvNBcQTrxkrPj0pZ3YTEd7vtJJw6b2jdNW3Ke97E7ZKR5mAvaEvK2kRP0FXx
TW+C99Q0qpxrayIGW4a5T68uxNnc4dcbR93gDi9BmnQE+4LHCOqo3I+lbBHeCAdH48z9FjeVHbQs
JL53Roy1CPrU85WqgoTjMr0inVndsce39chysqNIuDItc304BSDAhEpm+3RIjHlEdZZHrinvsU8d
6PGGbRljJ3ri18G2MMQK7t0kVhC0Gy+srz+iIRtpXGX3RtDB2SfucXPIm1V2n2Z3S/tn0VXiLlkg
8ZB8aWXJWDO1U+UWEsYoPpFA73snm8EgUAv/Tvzg5xiQP2aWzO4lzm2e91RJzq8vVF2RUN0v8AdR
OjmYpKan/ZCxFHqTbhuOMUezQZMAMxKcC/A9n6/WIEav1l5zlVUECX0xPLjfnqlFcaaSJs248vgL
JctiUn3JjB2e/9JGASWUQ/udrwF0KgvrDrqtgK6rLmPzmDsirjLuKtq/pfG2CIDZALkPMzZfpOYY
vvV8fQFvbuaj8RDu8tnOZ5KuY1ATzivcLLs243eYboltp47+HcrKFRclAwfhbTFxgab8tKnAwqPT
+tv8XI01g7bK2gY0PBenTaEHCDj/Nh5WsWSeIL/1EbJhr+ZGJG8BEQzGmG6k8DWN0u/4JH8/J1VU
iXcIjAIHnYOM8/tXv7G14z9UEdKNiP3qQq+rQA+niYSF3xj6Aj5XAugv6qR8O1gCfevgRlrwRIDM
3RdP5znZ7Pi2zuSbftDywFY7oJ8OhnqCPauAw/+ZfCtxWTFiyr1dR3XYisGDmnvgIgRfFCBRhVwh
QGBhR6mZJlSz5tIXmePkwJivcqG7Uy0EYTcWCNnP2aQwHN/X+/aPm8d3z41DuuSHnQgQS4eiYmE9
K2Y/ZrmyiyMTezZ9tHTzGFg+4dS5Dh6+8cI/f/X+12BDGxB4uCvkcA1zG0lDKrVG241KSrADmc9V
eXTrVXlOKixKgkt383qAGhBWd8aDm2O/8KXn0bKvIlg2C/Ik361RQgXYFBhoIrKIZqojmRzmwxO/
sRv3uQtQQ5V2m9nj+ZbA1WnxvsOXDvGel9vL/K34rZX4FTKrudIysS7sz5vDANgEOW+Eep0MQyTp
mDimaqpF1oYAa/B3lRq6iuki94iiGyDW0Wzranf0AlQkKBazUYsGBkXe7rikgbaWgh+jGtwoyNIo
pR4hBbS0Rl2TRt6dof5Qsps7u+aWCDjWjjtjMwXrLFpkK5ogx2gHlBehv0JO2VGIy69Nc/W5u3+0
Wu+IkoiGou5/qfuqmeqplikSKeIrbcDLN27K81pw7Oof5EB0JLe8sbpHHxRxbGrk7LREme7dUiH3
ZcTuB2DZxnztQUFpku21SfDLUPpF417wz4xQF7hICtdrb6knu5DuHcu8t0buRxHREbhe6dEK8YD2
pxlbnKOqF/zsJHCut1I55hcGZ6oerYHSDd1+ZdLi58e1RsCLNFg7OiY2nIDCLPIRQB5C3nkGJdE1
PMW6RrPEzdzIIgymD8EOUExHdeLpvtMU5OCA/vm5O7eWs7Gkj88RI9lxSk4nekejWtN6mMV2FtAc
NHJj8eG1THUsauMZEE0qqzDrvNnkXb9dlJnsduvgcsT8e7/xdfkj84f+WovGqnPOFRfjjaF9LnhP
EhEyO440A5kIYSzQ9s3NGV2O3EJ+z1Qs5tYJEkcQ1DCGMvvwWdAGZO0CH3Dm/Z37Mkyv+6OV5/Ix
dAfZ3VuUuri+We39S9JLVmAPwpSu3EY3c7se6YOnF1BunfbsQp7JY94TwfeyLabBigCPrcL4HZKd
UnTry8HP7zquVCjms4yzTuY9U1o/Edw7n81Q6fxIhy242ZvcH318b1sNDgxT0NDjO1X3KrLUop3C
0oHz7QtNkb+S9YYl4lRaik2UxFWsjhZVqVv7YoG51sWpPPHDs5fmmnmNQgbbd0T0Dau5cNPnGTiw
NSk3i6RofuOscgDkN9SVGF9Tnz4Am6Jl/1YvAdUGfhdf1vDCl2jKMp4od2SvZzVodGGQrRj1oxQt
fZI8vAe8/jqO0OWRtjxfno3S/l3ZrBAmHex15EUeYgvi2y9N6l0oaFEs+3Sjuv5meq0W2MQprfbB
jVuuMV9EI7xVT8rDqHKOhn3QLJCd0J/jHxmS86QehqlNwb4clLAo7UryuixpKYWoWrY39CfmZM2n
K5CKk31erIxI8SoIxr4nbHQtRKXD9/xrc/rGG7girWa54I9JLAsv7kvcsu1wJEWgL5k6eHZj6QPj
WUzq0TOHD3hrc+vk3rytZUzO+hUAKv33mf0DaF0QG0q57h6+I9gWlyGSN5AABAwHW+4/3XBvJrMX
eFHQdCgULfbyhToy5V30Gih+WT0Wso7aANv7JBKp+tH0VEEqRl/rOzkCvjDo6iqBEP1Hln6bfIY8
qW1BDXbO8tMTy1CeY9iWim4YJe7x0ZF+LVYJzWraSmHuaI7hN7AGGGEpnWJa7S6/rPhPJa+zY8PO
ip7YzjOmfoVwsvGTgPaSh8l69rvMYT/NDyrbo0X6n8akJyAUe1zXcmbfbbuKjk9lwvYt5z2viDlN
gekGKhOW9q2SHxxXuEt8s+mwm1GA9zJCnE3dhDwwlJQ1X/ZAlFVHl2Wbf9vS2k0jRCGLhWgQNlp2
vA3YTNl9pa5DOum6KU4UZTysoppFhUsBHBJDjS8QiKSc+vhMaOGUCesqjxoeGlFcpf6tGqzJmlq4
/YLd/H0ThcEHG3k6Xonx7aWbCIIVbqctqazgQs4biWaoRqr9UoaH2sP+QNWHzHntjiCGAR1lII2e
wpZt1EJeRROl6ASmeugiSAA/gZGHt+7r7YRMZCyB37TtfT/YdjCtQQYYFD0r+xmoM91oU08EusdH
NQE8ejjAqV6YsjY7kwaOa/lyOIubYmkEBnJL4/4i87buQFdDUxHTw96sYqvH/GdOlYJT/+vBLeMW
Cufq4/zhUaYEPiq3tmACfU72XAaJ0g2qJLB1+xDc3ZwtV6jXxUhYSnn8GOJeiWtayRppBqe3s1Yp
hPkd4gUT69suP+Y5LCAr0DfVdrm3M86gWaYlCu9cF4LB4pLOo4E0aaMWmbZn1NFHOLOIhBmdBlIH
CvNh2OSXo8wzZsNkGGDR6W5LTolAE0tMTOVHaB2RWOSB9iMj5/4dXPf5Z/aaWiW8bg7nYGaBwO/R
xnSWxyD7ak4uu181qtsvH/eODinV9EVOo8bPhXWdRyCVOxbB45Qh31PYxBPxQu/tKskamEbbNs4y
Jbzmc4hInPlrbvruAgfDNBfZnHe4NmgEAvHn2P2Oo/owWsyyUK4mTiNvYHue1gq8AObM0LnUD2Gh
j3k8YcpI/cqCkaY/aLlOKL6NrR34vEOfHfRLrFQ01KsdH8XnblQXx8AliPx2vtklm9vqU6JfnL4F
0TJ8U3weQuPJLq7hdVz3pE0xfoLgdLpLJTkZ4j4WhTTqfJt1HPUv/IJ1pTUzqKdzppSW75JRz9yD
Pl3QhYCvh02gRHOzudg7cd130ygwp/adXBTE+jW07BqkDXgdM7AqLGKwwjj3HHS7fMrrPzuoNUL+
HL81PIWOJRfGVa88ueZvqN2Z6pa5H4jJCzFvqEKtsvacWByZxhnfkdZWTk3I1pnoTV4JSMr7LqWn
6m2rptfYJc05BicpRv063m3LtFabTbvKnqyzNccxU8h9NfcknzDD6zmShUXpK5Tsp5FLpxtEd/Ix
NscnNTFtyQlTUQzfT8IgjJkkTIpnRrSQWSnevDeBYOQOuew55AS1bp7KCe0jZ3HehiWjGFsjObzM
CwBVt9hNKVHYpSSAguIgcLaVM9rZxSKSXpMIBos3eSacbEsQAwT4hUgLN/+WZD1QAqCjMPlYwy7e
nUq2xRgsiVGsMeRnQRiMOd7ccLaJ+pf+ybzIe6JFpO4JK3TLUGIjuiWPhdqooUscWX6kJ9pehbPZ
j4ShDEAfrUXfgPjCKo0eZjAtz7ZnyZYVyIeL0KgYSIRyz7tFXj4craGCavenhL2A9fSwI34qfrp2
XLdgRx6gfAEnjPfsW1vfgRWlX0NBi7RoAojbERDiZStMZXGUIEepIDHepIfzSuPBXMJFkM6RIi2J
uge8WZ/ovVLtLrb0OoAQ2mha4tHtH0JOSOLdcMi8d6DLpN2X+o01sKlrqoxJypTx2xRwUhIui5xe
vZQYj4HhGC3qrjihV4q+FhhKj7xkEfQqW41ViHyOBHRG84+I54+lYK4hB7/eLtQgCkYI1HVYShes
tz3cWTCaVoGHrEfqVfLXBAlZ8R4QbluuhTm/NeVsZLHWUZoL9IGk62fx0Q6BcAeEq+r1AndCNeWX
3Thw5HP7ONnkceQQrFc4tTxI/2sau1ouwZwjyvRgxVO64drsBTmBO4p/gulukR1tam3ZAwhec89V
G+s0e8ZrqsseI/96gyGVyjbgLdjkn9TiTMRbPaTozPjIwnWddcRBVr7xi7kEK+dX3oUxrOEWbcn9
ITPzIjR9i5roUQmP4AuICMiobplcZM0qk/4DeX5PfCC4INF2+89qKocoQpGgz52DK1hQluc/hza1
cFIbM3nYUjGhvE/zcS5H0L22kIoKDIdJ0w0Fi/U/9c4aGIGx4nU3ssAxGZIDp3SsCbjxW87PnBe8
MdqA97I1xBR/VIFWFdzoa8NEGEQiDa5kFUWbjnzDhs/5c3q8lNJSWP7GzuqNysXPUNS+vsviD0Ee
ZIFtkI/xF5fV4qZ9LBOXPrkj4CFmfOpQE3Cv64b4mr9vOst/aff7d9ZZ5XtSKX0ocxAnfjRufOLH
mYlqLI3MS5HI/NUR1QlFE6MRx85wnNhKOLvvbId2cqZtbFe7RfuQbvAem5wDF3zna+Vvrjit90fb
vGNJ8iXcY5r124PcTxVrbD5lCRB3ws+gz0+Qcpcobqd/9XBtIyqKPy3PCX+NlYII63roicXTWR7o
pLftCCiK1V3JDTgMwkyB100yp4V6CuSDevq0cuGRJpz/oGk+s2QjX+FSBk9eXylZoQwTCUla+bqT
vlKbBmQUl7ApjkQEyFU+9GECEHxv7KOEwiG5g7hIugARK4yylWc8NI12oM5kjnGoqity2nA1bnOi
E5VCj7K/Q83YOVzIddf1N6O/Yd8QvLseG4/EE3TC7gHCArQsK39beKLfhEijJJvdCyPb4E9QOqjp
A+qiT7hWNYUhdlvrIP7mdy/WM19Wtpy706SEhQ9Xml1izGZmDdE3vb+epjqSB+HVm2DSchEorLVq
CbaDU71R3cosEFLBGvRbT9/K6tz4ITE3ijo3EnyAJdaKHkNko13lcm/ddKhpeS6z0G3neS4kd1Ja
xCcxBBdygnAmsB5p/5aL1ky3NxaBjiEHRheP5z9syJCi3wV2ltrlNC1KL8FAyVrrF+liyFYSyfGH
iv6Si3Gu08eEAkG/3y9wG8nQ85y+jd/1/t7ZdlC6Q6ccA5CEI2HDNmNBT6gV0uDevf6MAQRT3TWm
ttF+ho8voQ8nHzURbQ1zVOELbcpmrxfclF6Ubzn9un9MMLF82+XoeSA7jDAbo1cXm3mc82BoYtqB
DLHseTA3J0tkcKBnS50te90yTZsu8KbarI+FDu7sGhIWQdyYw6vN+j0uztgRjq6c+P5C3HCbvkh6
B+iWPYV8g5YdOpJTtd2c4kU6e9fUrHwXuoKcrxfoFzOnopH8bXbO9Bg/2Esk2n+R0OL8kL419XbN
BxzQcg72bH0I93KF09+sFxhqNH08VRloZpSGNx9PZB4iKEegPatqOmp8NhN+DfM3ELQbhkvveJAE
AwW5PgahPcm+MlfHAg3wo4hkgSfefxrIpxPEg5BQl/+np1SlrYxVO7KMkekBYLrFZo2d7ImL8/sn
0RXmyTk6heQpXmue0unGA5zIl7XnV+zTqd5XdnYpOpAuozro8QDDH+SxqxUFGVsxFyvLMXbJh0af
JXhnPSgTbHFm83qAGIntJuK0kOKVLc8D4o0fl2zLX/cZHr+2ZB0PNLFAiuggH2ItHuSAQH8KrtB/
qU/KRUKecQ1iY3nBwNc4N4xvJZ14ybm4riRCPipo9+HiLte4NSOMahnhVTV0P6XxwgYVe116Fk1+
8QafMHTi5AKULhlwYjIvUmPG58O10M2kIjBZ57PAJ2ZkUUSKMvtOQPidTRuZQzY3/FoZMuJxcWWg
IVwUW8Rp1xbUe0WeWsB6DdSMJs00g3Hsbz41s06UToYVQffezYS+iufRmUNHdsa4jcG3CJUNpkq2
cMVHFni149NBjr7vQlul6mwov9Q9jNkC2Bdsco0L9WIgbdJ13djqNp2c9qmpPF7mv99t6MIqKtZm
GgcE1dupTzeSpC6G92vhLSbjtVtMI5yICKHPekHxQdCLxthvzDf/WHISKdiFBb8vzkOZpzeJZl9V
SWGRfIlzxg572VCCnx5dOJFFTFm8+45obbd2LL141L25W9Kb9ir/PFLlc2fPJroptq1G0gfvMrON
zB/uwaK4nXpDUagprul/8ikCLOUIOiKfg7BzC4LiDQVcAvPlaXQX25ApSdrBRd3V9ocwCP5Dzmgj
0xyaD+zwt5jMMKFDDYM4Prm0gCZv7lsY54S4Oc5OEJYa4vYdEiekgf3dbOCvvlMmYHhiXqHhx6gx
jJa5vdOd/1xpT67jVSHDk8DpKuqNd9uQfpCTDZ7zf4Y0Qtg6afPnTwxBpcbdasykUeFIUQa1zA7c
ak/fg1FpYo9UcBs77rtTH9vqBIDd520ZO0NJhmPQW47SVlLP0VuTxqluXaWYQTTyt2b4Au3E0ztY
c5afjTK392/KFpGRZFhP0lGxDDPa1DwgdwpKbDhNC7WXbj2QkZXeDfD+ARqWd9ew1n03eB10WwcU
in4G4HbWgjMRUK04jOcwcvA1NOI/qp++a1X9EQ0vq97Vp5hqw/7tsxNVcq9+Wez6Vb/pwIINQmN4
gCMgwP903vGWTB5qcC4Ygw/LDJOKxvZPW4E4QgVDl5thXPIwD0Nok5GVLBUskHp/vD3BacayxQ4/
mAHXJF5ZIYwjY77L+wtha+7YaTMek1vWqkMRyLgJFWp2yFj+osQdwXKPW3ibdP+JdFx2JLTa9o/0
NgB7j5NgZzCAj4ocUoloOQtqUMQ6Wh8oJo7bZ9fyArfjIFj1HbcOPr7YGrSknvstIGybPCWPzJFe
+UiVwEaTV7bUK5c0YcEAZTWhFrMuf4dyGsGI9n4C4pj3PvqENkHl8bex045UC+Xh2tUzgbWLq27w
Z30HAhG9RQgv1f4S6V1nNhFEhsBfWcC6RZhisvX76n97ccdBRRvF33YUBQCU+X2HLvYPj49E4g+3
bnBYaNEmNLEj3phq5vZ7nwPheU32SSUlhqfN3QGc+ReUUXdFDGhk7JjZjGMu1W47TdNHiW9Cg3IF
1QcIz/70Wg5ZRfHjv0BIg6FdNeC+3VJQaJJaPxOeXkYH2KcFPiUaKapAzH+hUemsuQ7oA0MMjs0N
f4f29sHfdHF9iWEr6nOrI6axbE/1zjZimYtKtd9sJuo4e2EYaEzozcdHUSmJF7+f0wUJKcWs5fBP
/pYp9IZdC3U6YdZeKToztv7fYcFnv0MJrVYLVQ91ICc+HTFNMpN90AVoS4HJCqQGqMhOCP+8ydWj
iY3f4ITLCSX3Z3LEn3+OWLDXE7QIWxIg6HUQA3/+2Y5sHgmFVl6HNISZ0IE7bTDExzyHfJg8yJHN
+rfzJW3shW7O9JZvH/gVoFlXfInRG3+3TcMYaV1sRucWayNapOUxu3Vkkta81sntNP25TeQ3JMh4
/85o2Cg0ubwmlQW8t7yukBtYHHr2hv9u3LrajrJB6PPaJq/emptqljzM5Ht5WXY0huhHZx+IZZ2r
NSftRKKATdzx4e0sK1V56sOcYy6WGqCTpuX2ABAl3c8QLhZ1FUX6qzTpGk9r/T7LFBuyBZs1Q3CX
oEZcbtnmyF50Y182yVDOliLqEmHRFTQYjjK2iOx9EYq/L0Vx3mzKVmJeOMGbd5GxKkqq1leFmek1
iH68zgb0gt/JkReTWL8dL4tY5x/IeCb5zyuaKR3uVPym3fZiKEPWZuvq3qxX7EV9xHDFNIYHJJ4C
FyuTZ1Qoos2ToHimXRf9LUYIZxGH3JCXuP0K0twbIv19Su1pb2197RWLbBZ8Ua/lNDZC2+reLRr1
X6UNKoGNPGYRzIw7p6at3s72nB9MgRlmBWpEk8aYdy00+FtwoCWMGhKTlfb55NkPET0yq3TZg30f
BWUNbeT+fGkHkN6r2xCaoREXSwmnjShJsaAToPhXSdaCfd3I3iAMkI0XaUB9O/cqGE4uH5ikSNMX
QgPDBnYNj2eE560BO/C6bAK8htVNUCZjMMOv5kWd3ge+IddtTP9cEeFK0IBde3B0GCp+LJtU+XtS
x+CGujSsRS9o3DRXSaJAQi+ocuUBiE79sWOIMgKf0D8lUcatEiif8aFw4JMVOrrPOLmnYXMzJWGo
+ZGAFS5LL/oncOP7XGOZLDF6v0PTo8HHSitfe3MLHuKYTxvNzOK/1toyz74tAse0QGFJ3Cfl7GNh
X1AJXJQEETHqGCTZpEWdyUrxDfsqAkYNID0jpgn1awQ/CSm2bQwDY2p7LhPYpAQs3XBulXO0grzo
IMggzOjJMGbZE82nCanTLJ9T+OaASs10Tiv7ypHygJXFY8FenmrtrJ1X+5FFMpnwp7QGlYPVqdmu
ebHhg3KmDqNkrIu4r8PVqa3gm8QcaZBu6jpYz5zxKaBbunO4rywck1kAeQFhq7y++ufTATAHq9a+
MXabmdf6f7Nyp6YekxBeZTtECjGC/6ZZhjEx4otaUMtPRelAP0QkUcol5+8yYgmQ1h62+0TQ6krO
PxeXjMzobAmLaD9AyXi9yrxi5sZupZNgLB9BjnKAOZb93Ava2mklgG4SA+eD6tNhTPAe0MWnYHfS
xj5YM06t+Ttn5b273tP0zjeOHhi0zlViNu9cESWfYhC8VRhmZMnX6W963UqdZCdPM7ldNQUTWJYa
bL0nA4VKS0pEJywTgviljD+b6LBmRkQjK9OuelwVDjVv3lSM8CeJjY1K2M181t7bqt1bG/1X68fR
hx23L8sfb3syPZePzBxArK9+PfSB59ik9VlUHXBWVvNDt9ueMBIpEqEdq63iWtBOcbKVNXEircQB
T0NVogJKxWdGTzBMLj0xx07h+0iNaGel5+gESY3vQBzB8IdnuzBxc+1VprbNReEXpyaFK8ezPNHz
yB6gxfd9iixFTJK4uM6CmPAH8G2DLPzhhNkOI1xbPfSs4mSwzABkr11jUKEf3ch6tmS9MA4+Ozet
QfgZpLowx0yJ2FIAyrQf/I2TBZvy5StJEIxz6LIZo3yDuQToyZpzMQMNyPcjxcccaY5d/VnKjHMA
+UHgqO1Cwz8feTO7EvS8lKOAosHRlFM6ZkqqkzCxr8JdjbFNWPNdh69rkxFf4WzJqBU1R3TA8fSy
VAqe+xaCfJwPXuyPmHsNNlFnLi3/00AofI095Dnw6UxQjA54oW2+gHD9NqvjriOJ7KdGzhfG3Ceg
yrd8sjTtQXSHg3TXr5dwclhbLJG1P6iaxZiGbfvS/X46RLxnt4+tZtoULol9Qp8Dz9Kv1wcfvps7
gMJndqJmcn9LvVNI8Zn7ZmjLXyQ9+Y3M/X8RsaNgJ2zm5iwmD6DBIdo2skjnhAOKZeUgNMPq4lF4
TrPG2cC00KeiBXIKJNQTPxYxtLhsDnDqo8+I/Q6NGLn+lCq4fwShByCatPN+Fbovu27d2DhmEK7r
cafAEUVpnDz04djl/zZa9F+BxL/q0uzUOwBFVa/hLyzKf3V/hmHR5Il4S4dYVJkGA5RqNH2HzYXw
W7aXk9OtYfgkybMDFpiciP50qxzrpl31BTvDcFyyFnSPzGIkQxXkoS7rqXT9ZaNDU/ULF4dpgygG
tnLxrVf7odi60ffcz3QuyFgR8Wi+svV/QzcGDa2V8kUQeespyf09yM9oD271DkvBWCwi8x6iwJ1Q
QcfoVJHM/HC40MXNdD+Hjn7/OYMgGG5JuVkBS/03JzCuZLm9e7rKD7puWogRI1jLdPmjGwAaPMM+
TocXLlxrHHqmKpAOvuIGUePbVlqxo4Fx38ZIca12XSozUvH889FG40MtScklrSe6vgNY9dI05fg4
eRz/KehN13SA/5T9WFZNABoJCDz5sXEXLT3l8ArjQoxmo9ZFCA7GOp5IGRQiwLGV+ykPv6RkTwl7
EoFHBFB0PTR8XsMz582Is7Pd6tEALMko4NvDTeQSioTAAn2T1lqsD7Bb+VPD7AwyuLk9eGH4c/Zb
O1AxrzMcPo2g4nIBhEFbAeRPRnoMnGuEQ7OBIdJwgQtP8DCVuh1yHWiXfg0GhOSbxjtpEdUY+xP6
sj0Lvyb0sQbFw7iLx6X5aDsrHI9y/34kQCvBvXl6vNt9qIEnMCtzqyU5wCeT8TM0tarDQrsL1t0d
FHQP/wV3PF3DPBzJ7zJ5o3kw6T8SP6LQgomy2q8vtYdaVRFzU1oBhsfaKe5uIeGib3gwDLCWe4Tz
tYXKgAgOlGDJ1TH/u7501We39wBFcRKPFoZpHWo3ws6kvfk0NYewNEXeiQR9EUcgPobeWrEPmhbf
XVxNNSqCj32OIuTFFXAI2ULbQ0z3MX9rXWu1XaMFw0ys4AcJ8+ALiviIl24UHGBH092W6MvRmcdP
NrWxT0EMCbGZJr8EFyPciceqeY+mJiPdw7JGsepVxd4AEdE85PYiHLbHy1swAGiPcFtRaV0w2h63
lU1GFzyNtKUCKY/kQkGou8joSTljd09COLV0pvK+jQ/tfD6USl9P49YPCxznyggTPV7wRxMtJxt3
VzQQofvJXIJZEFDbHOGpFH+cOJcgE7yfNulEPUFAsyVgNTW2F2fjZDELS3EdRXrDKStC68MkPilj
I9QEKjkC1lE2cBEl9RvFwHaXhdtfBRiJt0jaFD6FX8g4aUr8YdMbJKFsQyH2H/11iWwe6XDHWWbW
GXDxylXdlrHyThuWSPbBTfZk8h1B/DeNlen+LEGZWNmxyQtSplYK7TDSC3ErUABsQ83XSio+DRcl
19d2ECDydB1oHgmYDyWbBFFQ6iIiUMHcW0CKwJukwSXuK04GIkqVo/5QbnDhVdiKWQZaRn/9bkLK
uK7EuvrUW1hV8Tx2irAVAKgGJxJqlt2v9xJ/jnRvB2QHkZ+olhrqPVYXpKHbFvQJd3NaqVgq+zdR
h/D5zlvm23CEDU9QWz36lUhpDMdS2XauQOO1vSiKVWkJcM7O+6ssyUqthLve98l1uqQTvNuz0Z+w
VDUWsYWX4bj1PlzaP+htCnbDe0FKTlcz3Z+Ohic1fH9FwFxXmwxjS3m/MFjyICv/rCYJrnE+eZtG
KaDrpePSHuXzpIEz3pkKeTp+OhU7oyXRUT5MIgwlAxI0R2qHdeMrQIIifs9vdOPUnjJq0eZT85Y1
vMnekQJxZYbnIAmpuRYr2MgftBmQD+L6HdeFqv5n2HNM4fOr5Dco8y5Xfi+q0Vz4UNEViM/1EeZb
TiHOZ96mlfaQibZOCVoVVpi5kxU/f8YPsrcbyKAaQJvDXWWxDPmSwgaQoN/XZThJRusn/T2IQ/t0
PqzrQw7O+dI+vrjyDT7Sh4rXaI4Ke7+lyFdee/zMaZj4EAiSMYEDTu1wjwjbuHkN646mDS2BWLJP
kg78z0mNcsjAGGCX9JxPPunghh5kKjwm3TowmnXdH9TCd+2ndTFXYDlxYWnd6rznKGyxpuVfUQBi
4ste8p+Lx/14+bzQLnLpa0SOvqvAGq/U5gZU06fxkveK2RFAJpeHOBuEIRkkSfVVDc60N1f55r7v
+16ciIuNR/8Ta2Y3Y2zvOQr+Ev/Ei3itcDAHF/uwHF6EY1UFvh6Rbyk2LNFiu1FlWlBGQX/caqyW
FGFOgx+AQod77ugBv0czX2q/8hDuQji1wGxj8qZJgcnBHYnhnriQZHC1VsPH10/morZHqFenrriq
A6Vc7VtQ1RsMtpIhYWSeVe978qXNBE8SUid40jSAG4CNiMB7jZNTVxPcGDfuMaW0QgAuojkLrBs3
dAikOMSBcoIfkxJMFNqEUR5kGLgQ9A5cDcL9xuHGeMedT4b7zG1L7WkCBuC8tGNyKTCfN1WxNFXD
ffow5eMh/+dbLgX6DsOMUKGr85yJV8sbUtj6OXbCuGojVuQkAsvMNXHg2OD2YIKVDkAtEbFZIDCD
cjY4RO1xJiKRq1o5rvhJvy4dJBpheADUcUglFwGIS2lkplzd1vsxK1OHceMeMGTjJOxy1tPytYDU
t+Mot2buIXaUH563TiPe0tZOvTO/GD4t7sNlYSb/ZyJDwDcuCEgSbiYLQ3Om8F7PSoMc1++PS9Iy
BvSFIWe9r6UBAGA3LOr/qyDj6gb5FxBvjjBFTsJe3qgdet4YktMbqVBxuBLZC7MNKijg97vVv9Wd
TTu85pJzPEBzNPP96FoLLWb/71uqhIfIRnnCbLcL/ZRfUt2y90b+7dHRCtucKw6ZXx1Ob4KHrSXn
PiH7cuq4KRr0azBpTj7RYS1BYkthebDw0KrrRyoyvMwyVyaKmRVp5bcJxAToL54S6ewRp6FAE6A+
tCApjn6HAV1lOyjmKSL/r12rh+WkdK7RABcVq3mk9Q1OaPeTt+HNbT7nFh4IQXCpTAQrUBac1+HL
nZkylMfIMS4WqdL+Sypq0WY03LDY8NF7tKW1nTeRZXqD5SpipvPLOiHPNOHoX+SbDOyorXFmYh9T
E/O3nocDNpim0XF/5UPdZ0YTB3P2t8SlcIejaMP6XyXx+xQOBJRjII7LsnXYudAuiCDZ6IT1lQbN
mo5Lebil5HNO967i6Vi07KZLzl9xqAAB+QNy9JUwFtRXeeWW0v8funuQhj8l3ksneluKlsld2VSK
bAnZAPFjKOTtG9UGO3rTidvWAQ1DgnpMrXa+y3ccW1kPGaApyK6ev+O0eyCifyKze9zbx0HzccSp
3AWNAvSF5J3bFYqaHXPyxxRh/aYU/IwKGSNjBUGps5UgmWmEb3/BaBxYW9MCRmS66yMW6+fc8Pek
cAiSs749aKjtF/3GbXW4KHeNnEJZ75lfXrwiYpnLvwAc6VPsWZ+NnkcJJXhlfw0E3qAoVEEHFSMT
me9Up7O8phx+ZNZ8jRgstk+XoAzqq76H5QaBDxLphElcAICyhoLXMWqaOXnxDaEO0/8FyEc2U/v4
21kGr90hvClDY/miPlNA6BHS9QSgzy9YlVFyZvDshhTsV7AYOGwIc4lb4CX2oru8+kEZUiFujAux
ipiZd2nJF+gOjbXnsO9fPBcg6KNSoCu5d99QZdPpUxmwCaD1oClwjzK0vHgm+FWri80nxde7qWd3
AqNDb430DN6wbx+dNHaemtAWQu0q3hBt7nwlxFcG9dbu7ll4TLczTl4krSMg1fqE7s2iizVOdrA4
YT8w+bxFRo28c0sbZIzpd/4EBnv2YOQUl3ngoGvP/3ggXYodITt+NAV4ciwcsVa5EBLhcxvPewCF
ToAeh16vNuCr6mFM5G46WVQbMtdSnKAPHgCRYerFPasbfbHdLHGyKw3XJzCtVkcOjbTdj48H4PFj
c4fuMkLTe0WAfXLif6Mi6QiPvQS5DPpWe2sNLUO5mLJdrVkUdNXs9ysykc/3e3HR6dbb2ciSPiqf
MoQo4a/C63opDOYNS8t0yGz7DLmAGYFSWpoQBxkLvaalxZEg94p6nSglvEucB1BsKVTK5pg67u8v
uFV4AoiA5gmZA08BSV01RtmC8xk1uW0BtERmoDEz0R60gk7eRTEtoq3K2dAH04XlY121+BEZBTth
p0uvX+9GJHMKA8bmxikSXt/G5x1kldhMYF+hc9MjKiJ34GK3b7K0Q8FrGKQ9xrliAg+6XrJ9PYpe
9o2pfpK4fPGzJgpLp91jGdk8Gad5k6RkpVN0ZVl0cHsS9MkHOlZqPekyLZKXXvk3uwyOE9wCsC7B
ReHRFRsgl0KQLckCNW/0fCM3Wr2SRWdRTz1V3njCAnVZBa9vgEvQawC5mBWGNEN5b+ZMoBd+1TzZ
PwIdkT0HhqF0ZGQ8QOuVnRPScG+H+c5p6sUz6F9vMZdLAH0kM9ga3DYZZlLpifhnqn6z5/jY3f5R
E9jm2Z1x4gCXuJMOBZQvrI4kEwox8ogwaZcCXxsI/0wELm+977+MlnpqfJ57ct6VuSKj3buDTfHj
o+VcZuSUuJ57jwPRnXe8WZPzHEH3xinY00CUTedYBm1Ezr1VsaQ0wwBPgCfIHQBvNsUpmSCTrq1y
iGuRGjpKjOFFf8G0yxXymqyw2eXuiKcTkZfcAoSKA8yCc+KzI9p0DoQGtmO9dtr7k9CjtBMpcjSF
SMOIcw6C4HNCVbeJYSb2HcoLBhsTXO6zQ4mBXvFIKvUIgJdZd3FQVsQNDfK7l+Ew8FUh3Ia3KDHa
F/D/PoN4HR7cLFB7+kb4xv/u8HTvhJlRLUZkmMUtEpRVS8j+fB4TjaztgEEmbmPeaaFmzyDPBiIQ
NZmETJQIlug8Zk3tMqQNbI8DW5IMoD9+NbRcdplQZhdDIoM50B589KI1GfW0RO5vjrpIFpaHHpW2
Ei4F35rmLWwb2xPqp3uaLziLeneodkzDMBZE/2MNnXg4KDJwMZvgCg5B5KKlm8ZgrQkvFFYyfOC5
oFCjq5178s9L88vZMUNbHPEprQ3CTHyWCJiUMer17LJUVehyDt0vD1KqDOA+mtVspw3sf1pBF4XN
oZUN7IslikVf5iUIhFDIXm+CjV7lYIis3RVQ444KnluhrAeYeG+YyJ+L4l6C1qdw2AZ79iG+lCfG
a41szBfHRJw5uhSZvKyIgrVU5etXveKLK/wDU9DeXn0u6SNx90c/j8n7bYrUniygLR6iRnokVheK
MBuShM39wICm1iQUaCX9ovo0XGEQGbozOTZWfes03QK9fGKYROfVXB0aEK2+uWFKh5VuFeh5ezp6
KFqRtFv46D98N2CE/9RSRDYlynneseV8u4KeMrrIfpZjxevVmAl76HwIWQGMzG91aThbGXkp7xXa
ho1r6duITH/UwMKbl1w6RaDXqZB58caZjx/eWB+hqSyOPxwjtX8NGrw4MeoKjoRRVr2KST7YYagA
cHDEKYB1XL4ysaUqD+iLGuD9cANsB8K9F9wL5wLLXpfdaFl1hDMdRAtrhqKA4VwUVVG3YMU4XMd7
G9nk8gAVfhxiyR2wAkdMOfU0CwJLXncSFWSOx5PF6icb4V55KR9fDCQfWdj6cMYO7M5/MaqBUFw1
I19WoFUgnFqD/0gM5F2PHs21nz8i0TCBxuIqS5VhCW6G+w+W6jjGoKbh12RTvsJN7x4IvWW6YD9s
iMcz2mdCzTUTO0UaqBXi5tRgxbchxNpqz3Q5SOw5oO8pdb5UVH+h/YwRmpdO/AyOT3E/pYk1Mbet
CGXejlcUfw4NReP6i9/5PZVYFUSgw1CionLzGFbrNjVwh1JeV5/1IdmKqzXIfu97HIakcT0xvW0d
wQJlc01GgUSeR7QuY29nL483d1dTjWsy1ie725JO0wTSMtJ64ZxQKmzTT+CYlWKnRpW/eaktDKW3
1mqVAbH13NVaWPrMDRx7i22ASbgcNojUkpWzPxJ+Y+xZ95/oNPYgDlMKl0AHkq67V6i2zlbzc89V
F3GH9YQnRycr3lIVpT5kLaCAmON05dmFTw2bQIKIozwtFFF/pR5dhE3jscD/LIDYrch2jd6rgBJJ
AWYcFtir0khLA8w3URLeUlj/WfBIQrVFYJMkMJO5SkFu4ul18iV8FCL2kAgKoCNdABVC8nmq3/9q
sGTWsMhfGuX245gkMsJoDSnjEyFesflf5V16FBIeUm7Mi5rcb1BSUaVe6Dqo2Eer+tiatcDP2D01
Nc0AtZBbj7h3R42zyAJL9SocfLcq2jutU4I6ypiD5IsfuZoN1bCMBdoXUJpM6UaL6DQlkQ33JJ4K
1m9oPVeYQApgo6MFdhJKL8yhfzmqNNCQaGN8kdD1Kpe58yL88Ej95bGKezdJlz8WGnm8u70PiKwI
SYe33+JPpwpbocR6G4UmKjGApwpd/LGsZJ5sAlnZuT781EQV/tzQY2yx48fLtRy6hCkK85X7eLqh
DZVoXl/OtxCJmk+F8V1gggh6IS3tn+k2VN92gs1vzfTyrpqo2/j6An3Fvjy67x5dHlrUU+2M3kM/
aTMyGd5bq3peb860b/Gl4XsINJQdpphuHR5llkVLWp7gcytJrgkZUWMY+bKE4WLapHtY+v0mep0/
Cu7CG29OplihAf9cDUjxFMFWS8YuFkkf0T6p2xIeeKkCUtB63aBWPRR67Rq2hwA7f+zUPSC92hj+
rIrzVDJeWHIPWBwR1K+bMP7WiWW9IrtI5zRGosxP9zlGfOgIeZLhnqA2uCcJWKxGKygN8A3UGRIf
VeIO/EwC8ZElZocvexeBbsaBLFogee2GPAvv7UOOGFzOEdVYFLsdbYXViRt3Npi+S2zmPyLeXdMz
xI18//RDbckV89EHioCK0HrCggj4x3/If34eCUq0DDUF1CpC9os1l4LYL/dIvRUDAqxn+RRHBUUi
A1dP132X+PaU31c9zau5YgB5kcyi816YFQ3kUlZDHdssH3zMWk8NRXEkMbq4akbcuq+yjaachXgH
Q8SRlVw7xmKqSr9kMoJGXHSyFxy3Af3lvnvQI0VZDwNPUtqaUiwyPdz4XHUOV/VhHU1SXdeSnjM0
ldanCPmpiYJt2TmYnKNEt7UfSvUJyn/sJkwdj2bQgPRzZvj4blgIVhe68TTJ3qXbF1OrN7xzY7qm
2PlTMN9KDdA1vSjkGvONDqUxNR0ff96PrXmozCAMB9WAAS3T/xgo6fIxC1qXmhl7uX/EL1/PKl4V
tMOo0TAH4DlJU0GjuC3KDaY3g1yW/xbGZT/pD6rgz/qCGD5uNzQCUgZzHf+n0bEhsvKu1pnVYP0+
KxN8e8irLQyjc01HeKIkMUyQKaKFija/qDqMSqYhC17+xtFMkHOfHwD1BePngQ8oCylPXdhBdrLv
nl7i49nx6/60o54N4A/zsNeucLfyQzsUssWE6V8SufzP+Bqd1XH4jwF2kaeC/ZGcO4MMr4K+lZEX
y94dEJfIlUcN1PQLpzQsmGHKtbT3vTGucZy5Ip8uSuvtcGcKUCMHqYbJCFseRNUPtsu26E0WsCSy
b8ueXiScWpCoxkAlCNKUjXPQbjcyJBhx3zFd19RKQ8Sn6nnNK2K8OMdX/5Uc0kjCFHYf9Ozd11tQ
xSXIyLhcldzom9rbM5gyrpKUq91VwNUhR0Wzoz3XIOWP/6dvNfJno86u4ML8CfSoOM0ub2uF4nlt
m8JMfA7eVh4kEmuuLdW8R8swvBfTAj3xnxaqm9SMKxeaD9psy1qNn2wLZ7g8v7etYFH41A48WY+A
raKhGqAZl5oTDyVlO6vsxldVBBndiUxfkTqpH3Te7ezkIdy0xMWK4xvM/Sp+QfcoXxCSP38jN8+5
YD1UQE3ZfEcAVQEF+/Bq1qktqwi/j4nHG/uva6KfcFPVOZZxmAcEWLWxNRv9wsbcTUrnHLJh/4jf
6Et7DhT0LhJ3eoEbTsJuaGJ1MPgn+vDG/F0cb1GNIqDVjhuS7pF3LDCtRCK6eo+aJrrhoPBPRIEN
qXF5lLCiV7+lTwRVcpiGRW0d/KCzUNiNoHaQmgGlLqkGZvfePTS5WXW5zf/S6BtaYKbonvn41JWx
uicVtOoNh/53ELE+/7rAH7MfO048QTpKAqNj/bVk89/UtlxN2635kPaSefC980Z4xMbDYBH+8X01
aMmRkqUZMk2jGQ108gOS/AarZQDzZhb2D/mVqG642pMPyln6hVreX8Q6QXzkiNBXceZ3Pp8PGGOZ
J2VtIhwEP5jULx6lftltwdzvgwaMdopF5R0t+sOVSCCAMJMgW6k0WxZBZF89fhy5cF7HAFLthVoo
Hp/xx8xP3j3yCS7hfjLeZFY0zE2ZjTDE6hQXxFUvaUda5MS2zMPfyzcyggDZBfaDteh3VgheAD+r
zRw3OzBsK7YRH6qf6pwsw9XG1luzP3lvOVTRf373EDVb9v9JOz6R4mjYTTys23uuiGypp5kw9lVK
BfYHCXKuldiTDor6F7M2FOjewDV9LZP1Dc/kjNrtZyIg6/wJ1YYxEpQxysXWqrHHN++xukSN6Ee+
wCqijg3gX92SZF5sW+nQ7A/ySM97M0ihr0SMyqjGzLl8i7d+TG8FSYAe89iZHU78rZ/vYgKSyx54
dPrCEmdWu4chz9gPlRgZ+SlZYuTledLX6fBiUiYspUPXIEn67O6qLvt7D7ihZ7SShrimo6bfRjey
ajQQC88UDvlbNsyGBgcFa9G2sABUa93pZlk/HZxJrkvJS2XDt4KdtJtKdLcfDp2gPfmBzzn68dYp
PQYMjBHn8ac1aDZXnIylrJ8+NVVqQLfezQaYJG6DF+LXtThr7kx3XMoLUcIZ7Alv+9vZonGCxfJJ
qoFfhuK7dMyUdTNR9QOqtqIRCkHlvKVGMf/+P1f5SFSVvoMol3kS4OgNqztVUef8GyxFcpXulNU3
It11tIpYqPr/pcIiz+v66TkGvr0miBTFHPVTK0NiWmYmRcbQw/2oe4SDs1JEkrjb4VpgpjOuruyM
T7M2lNKHGq5b+AsTTu7OJfe/F4AjPTm5Vje+mp+hOR4QDQJaUgultMvIJIsxDDwMChCxyvHQRDYf
J6+i0KkpGb+7VZMhbpL07QWMmpSOuonNtksVPQRwlF1kh/wxohzO9352Kk4WroylnI9GACPYekuG
bpqAsayYQ+hAesF6f291B1JrYFmyhTnxZgrWslEmdBMi+tC6NXkrJbPBW5+sDKiRFt9h/dCXiYuv
+fEtqAN4e5PSrVrXVNJYwESzjdRL/hdd/3TIiMzCCXIK2lBoFhqeufp9364/AjlD0L0rChRy8onN
l1cDKCGA2Shza+Bm1xq/hZqSdMENwLalN1PC/8vsujEOmR574jWhZmhsh15zW6veN2JlBJHBywl5
jmGoysmCr+VbLDdy9ueqaqIolCU96GBkw/VMzTCJXbcxaaAnljN22reSmKykI2Ht5WRUfRCx90r3
MkRWezglk4obkf7cZAzeS4wTCVZ8rA3GACz4yYPHja/F1yaqJDySbAfREQHn4SceSLdMilm8+i+8
rQAHSnmaz9PElytn6xiuX2oTUl/3sNEWGYChx6WAaECKlQbq/Pq7UzxzGSU3L0bD1ZoZ5CBSlnKk
9M+/uVXcKmC1UqbrYuosJ8g9FdLiL1g/jjw5XSyLwn2Cz6aOa7jEDQn4NG2dDvRSfPGVSLZlR0Jq
xPXLLvGoGkjk6qBetMmOiFtH1G8LIo7j6vNwZjjLqoRIv0nYn8R14mfT1WmpUTYOIESU4ycAW+3Q
rBbZCMpclAC9lK2iVhJj2Zezh2QgevX9o5gui0+snYbdff/3MNJir8PMUt+ic4OoVGCTG7iG8Eau
/Rs+S/bnnyy/g0yVqaKp4JFJqiI5Y2QKzj7PM+lLfS3gPXG3qXQTdb61UGXq+F5jE83UF31iz/Vm
tbOQw58oyCd9yTEs9p8L36X7uWtydQ1/gqZj5+CqU6KMhes02bSfJTLjzSsS7ecQ/aQ7FNvOrqUD
fMO8HoFYuJueVq40EfKS74eM8RdGfIvnoWu4cNxqfnyC6gMZRzpuYVmEbkO8U3tlZP7T73CRBVPb
wCVHcGj/TfQpYmBqjiE4Dre+97yAyk7gYtw1RRLw1egNVLsVlYNIyhH+I3xay8BvMd0nZ3HIWqBY
/vme7BvWn0rP9w5+Lvaim1dzyvQkqmZail0GDwnpD6ZAZvbBDomrazCNb9mI8OX4Qf/3H1IPKVIN
UmbEh+pj1MuNNZllKogpdMkAK57VDDqHjJhylCI2JkiBCnOQqf730dAao9udcJ5QjnXMhi9ijUlf
QjqA5y/S/Ly4g0ieEiy1DKir6lonLXWy217zQNyDVE5pUzxbHfMPU5uqJzKLOrTjxRaIpbusJbXT
CFKw6gCPnxxpARp5DydSi4smgZ+ZJOpuHHjGEnQ4xZr9bLptUBVEOUXWwz8luc625tr1Fb8VaA3u
QW91Fw0M1uJc/F4KivVh3c1fPSV2GM47U0oeoqAFuANTexzFWMNGR5vBJhWzi3iQXotblsrgIJQD
uJ7bLrfVd5nSq2UgZRCQVMS5QVJe1biFEoieBdNVgJQwDulYBDjae1DfaQo3BMIPn6ZB39zgSW5C
9jEKQ3DlJzfYs7Yl+vxzBecjOIch4deYA2dL65wosj9553y/QjdO/QV1Z7FJbGbd7xtFzCh+pyi0
2b057jz3rfRgPl36CaOPsmxr6AzgX/9jDZuUPP+Ovnx/vnMeQH5I9bxCtpjdvFO5I/ctiXrUSKwU
IaokA/ANXIdv84nrY9FraOf0RwtSNj94W6ugNRjNwqeZnjeeYwaLmrW1t+wKMi2uGI8mK1e6EznF
IJZI2TCsEKbfTd2IQO+uoczN1g34AkHZjzL/kwHjIvxEauOYnogyR5hajJWsxCDcl8yRs5vDrzbl
MZmsuUrBKS9n6uxhrPxRS5Uw3XER1ZKpKJn83DtFnpeadzXZN970dS5h+3QQjh+tdqFTFZLAzXeI
8Mnbv5AJoOn7EslvEAJkbdbB8cFpSCxJnVJgsqUSJwG7YsLqpaW0PXJy/HHgH8ZiYR2PXhRbgusW
le2MezXOO0J/GxZ0Shzqkm+qXi3309la+GMImwAPvP2oMGQH98LBoddX9L8ZNI6Gh/3WaLMnFUC4
OghKEe+90x+fEnQWrjyHcsFNov8vKtkFjGpq9XJVgllsYQIt2R5LpQg4X0tsyhUlDgT5iXKnijyd
jIVgFcipaEiVzNcak+eIMtzJ1YRAB+7nXyejf7RlrQnmQ4Xfuf+Nkia9VCFSxpZD/8+tffBXw8VZ
9KNOI1WyDZ+XMyTZ8U4dBiM7+Sx9CiMvLelwMB9lSaE5PkI4nuJU2jQwPVmJ9qmR0gJoh6I7QlI4
TDs/Ojzx3NT1H1/pziMdLwxnpZRnJs+3GoATtebjkRiYONcCif7GwsLwMnVx29vA9fh2k6/0yK90
KTGliOssq2OR3MJF3OZaR7ZPIh74yHXhWZbYh5cV+cKP7vUyFVGhUtBpjbXgcCwWvryfLQecwoG5
6G00ActWuF+K+nFk/52jZhTCAEj+lzqrzjRn4WRR0bkSOcSw/uUULJ5Qzgwa6MWi9vCx7joB4XKm
4E18PSSqe+miAUlmrw9Vd+MMnKpF60ISIuSXSLS9jiEp9vwHsT9v66EaIY8PhgLxrKW/+SEYszWZ
61fwrKHI5e3NPaVPXZveb3rtx0ZotqzPFk3hs7f+FuzpRISu3Bfc3j3/iqpDRGFaVyLG/IeTgOjU
bvD2788e5mYzF7IhB0+7bY+kHDBjTVxsHlRW8+dn3hJRXfdv8U85M02Co7f4/MIw+ZzFhM2eWTEo
iTFmMgo72N9R4fkCcg20whml4dtVLeM4dSCDeBzY0zEYx1RMkyvhDpq4gEkV2Pfi6pp2KW48S4hF
2Z8iuVqKuglRt3Gc7QIGsS+sw4uv7UumQfXmxsObq3pIO//8KEQoHwM3a3+OP+zvsl+CETJP0zq3
hDss94wre4EyYrf6VAhmSvFgLeZZ+qw/RXPuatD6Gm1j1M30V6nFAjzLOzQ2j8QUMPFqPuONvnsS
GXKjREOFok6MS3tUW54XBF+kvghCV5mwntnUaXPj1qjo773rPnD2nWWvuOhTiHNncMDuhk2iCHXu
liLU4duJcgY4cWdGFGFjPKUmMMKLm3c+YBUsIvahNARw4P6xEMt444RsDdRR7hSSr1mSXyGmFmho
pZVaB5wM+/oqq8ObC9VaOyUVC1Nzoop/B6Wyhc7bazvr7MxDXL3QZwgCt25XTjrQH7Ag5IXgIwu1
2xNtfUWWHevEJdsuP3EzA7TwGOO1op2892jNnmk/WC5IDKZqNjjaGSGE7g2z/U7gM1W1vR+sKtxO
7Fa8KfiudRu4Caj+cq0d/+h3GoPSnilGXNjd8zZEApLXY0YhoRKbhwu5AyJ/3XE3T2k64Bm9aG9B
WlEbmnJ8Of8V5C2QiSXWNO1IY20oIna1FhJpOsq5j4B5nhjvFuOV/8pTpgZdGmFIbbvJ1gYBqgh+
2KL/N6+3YqBnHzxuBU1V73RVfyLx+sfRcglFN11tVvEyC+uZqRc+Csu7en7NIxURT/gFIEqrcGc0
3n6bUvs0MKeJGbxYZa/alSkNSobryfWxbRju+cRq63Dc0VSVDZjqvbZg9/eneg3PlaJBsphy7eBZ
oNTeTYY8UDs/GpR+Q4zVUNTxrTcbs3qafE5QgtynCTJgkyL/j6PBYyoGK2oIv7aVdnH7QumyMguE
gEm161nqVt93K9w/d1cjwCHouApseilHtTKjFkOJRTTrdLeminG2ACoOG7G7EZl9AoKeeGF5sDkG
EXULg06EyZug8vEGIpXjVhIv673fkRVaTBFGLfP+Yfw28FjyK/Qk0omxDJaNCAFEreCCsRd6dcnD
6852c7xmEcip454GlYsEK7THiCgORfeUCpBS0ANNF1im3pCWTkaSxtPcXlWX76XBU138AX7Hdzwd
+wqlxQJitPsGh9yRHdtm1FzAcfjLD94bCFtya+LAsSuL24xzWxqo6XuG20fVXMztRGcRgSQuqAfc
C5hQ9/K/T+PjoDOekx/R2bIGO2y78UklzgFJ2YvT1L/ojiscueO6ypNgr8d625DMGHaOs1WxC/Sp
zrtRmZA3N1IbunHBWpOPbyI5dHSIpKm8VR3rlbmngfzfJXZNkMR21WGp4OOkJS3/nr0whPk/yfWB
vlb5RZYjMgvK4RyBUPGp+u6I3VWtpSw1P5jaRQHdp34E1cw3zu0EY2VMdrbkvOiNH/dflJn0atu/
mJd5P6EqLzukNS1Czm93fr1k2RWVYKXrMV2ok/fPqiaog4ognZqpVDkDY+N5/U/Q4sXMfYGfuCHN
UmmAl8j1zzKew7OGcwOqSC2pxwHl84mV4rPAJJqhCWX2jAdY85CmZ8PPu3OKm6Ysug8904rnx1yF
Lqx3YAveUWKLy//LV6fujJV5xtrqAparZs6gT9ON6L+OhiGsmJYcdAsQxBteavVJV2t5AjRM2+Pd
i0rLfZd4Ynfal3EVm0Mj4G8974xoovKjU2WBpj/Q89ZbVB26D2YMoxJDDGYsaCPB8/T9gnxwRUvU
VlKkL0VXv+mpch9hcVJp6uCSsbiZFqa8QwODMF+wVraKH7N6/Q9JKcNdxN1yiG4VsZM/HndOS/fS
YsYxaJfahFffwCVT3WPSCVnQrSqE1a7pjq8PkFkZSWWx3OsKT8KQerTz09hidE/GEr4131DQoD+j
612zW18vXMWBX2tghKr/vvDUHIVmdQG0R6MCm8Hd6Gjt2oANkLmYh4fa+pAcLm1Cp6odJhlpGX9I
NfBEw5XQ/eXXfWCWxvrx2IArxUf1QFU6oPSPLV6Kp+eETLWsdsaYq842E/39kSjCmIRw8iej92WF
/FGTdzE6of/pmKFwTi5c6UhPW7LJcz12WwUdUBKTzNu1RAKKeUlL37TQTw+Ky1I6UUq645S1S/3R
rwHSz6ya3B8QuCKC797GomQy+1SDQabza6j8GU9LVqv0TzllWMyGArwFLekuxBrcLZ0Bxv5ihssb
y0hJUlHx/jTab5GU8o3B6YmJcn5WT9W5JOH4e2AlLt70r0Wzv0QicS/2ocI21Yr6JH48yvR33urc
1LTae65QD2BR6/8cIwscpHrqlL51rMDxz/LS9j1jpTv71GqYFAx3ZWQB47q2Ww+YINGC2xK5jNA5
k+FYkvg96itKF/JVmzhFe1GuYBMFisu/Ql/o4puTOX5kUHyzLErjdJl1oiHnCkWaVp/7x45t9P8F
Lm/IsyxZwvyBR4d5o2x4fml5rD07H3kgiD8NPMNgaIvcH00/5Qmsqehv8DQgXTrHo71EDxo7NPpD
IyTYp2MttdDbMuAtOfwmQygEXm804cQNTOgDV3yefD/wgljxku49TkfU9uV3Q3ypc0zC7zgkfX3B
LmOqQIbysAjMpHKJLxGayD57SknX2FMY3sYe8o4qE+gBMVhSeJ5a9/NVYYnKanJscvGjLsgh9NeQ
xMi6IQQO6iFN6FZgmMVt1EcldsMDlhiEcxMxZxPFksIUdwiRnOJ3eBLDamk0tG8rtKlD8CnEoErB
S55ceXNs376eWXCu4DyCpbcm7B9t5x3EHvk32OS21bHmRCr/PBET+WqVdMvOOjm9WUuGHVrpT2Kh
+ThjM3zIa9f29cow4kXucglfHEtrC/zOHa/Ep2WzeX571AiEBl9nB6zke1wcyhk0ZwZCulCFj8XS
o0k0eWtMReEzKxyCa3dx0cBa1ZIkSgNQi18hlLr/r8CkZu540Gr0py6R6lNEu9WipQqWV/PMhWV+
O8qaHCE0hGmK/kgQHHRFycXfXqJiQXTvkjv2yS1QYUhxdlgUolfbsciZZidUNiHFVRSTbWaMiclh
O7WZOuzv3kxdWUgd8jnTL+gRRMhIuoqFvd5pwf605sOA+xwwILgjkjL/AMpOFsmDceouaTQn6NTr
8VnmRlA0rwYprxS3t5sk9Yoil7bNKkNfzHAuD3tAgvpQFbtxrlZQTJ+kh6tnT9bI/m+V3XNFUDC+
u/inwLs6UbXlJBiUgJ0l2+2dj0tneUjJF8fZZuTfpdLx61Y23054FQ/ocOzhPyOIjUnrvCqE1YpW
AUaOUjI4u0orNuHwCwGpa5XhaGZScQqxlljR3WpxY+sR5d0lJvsW6rKuKWNJnzsN6j72fGYXHt16
kQxvCZ340Y0ZyW+e9j5QwC4f65VzhIHnQWyFc33hGJOnpm8QSKubuZ5d/hI4SvEVMh7QWWBwdzeq
vZ4jjOAXvQnkKh6Xo3NRvxH5bLQuSFINaegshLocP/pB+T4tt5ry8I+NGyzJRdK77VQHHthsoIXG
AC6dmjlPqiU2GJktfpSJEqvL/MTMdYQL+fRoucxn/6gGpYoWVw/s4hWGb8mli9e2QYiubz84uH/E
JPjwnI9Krt1Tf/+VRFck7OPmAYjWIUCUDrCc841/UPcM1EtGBnHAuAJuAnpCkdv2f8PzMshKRuMu
vw8BUXtolQ8wfKC/xM5LuWDvPcld8Sf/EM8xUPZWqKoXV83r+Yh9bBkyaOQzkCBfA1Lxfegzl3vP
CiIUXDxN2xsQBBxrTEjLNIzdE+vGkeUyluQ2eW1BGU1BkR9YHTTzgFUtGtp7KVcYpExbHfyFKbfN
5GzrgLke4FGpZOk1Dgc9xUQUGbQwe+age11Si0L7LJfxWstGjoguACv+wLxdE4O2/EbxAg++v3Zo
PcDk6eRk+GpxmprpXTgNGafdVqA6zfvdjL9oOJA4D1skm2TyE8EBWab/RD6X+HaJXC1FBWF1ZHOP
MFBkBScmzjjHFKGlHHtFAzu67tUe9rfbk0DfPV/lYHyohMJvwISbcgWO50KpGzdtQd3mZJE9tCMw
cJiVH7Uo5E8E99uXIyob8xbketXCW1+QBC5P+bAn2AmfMxzsQjN2K9hbfQM6zePucHW7//YCChXh
HDT89Ijaen9cSAFWk/S0tNOw+5Zc4jpdEvMJstFmmJNEfYQWvNHYXRbiQFuzysdIOBA2BLNi4RI2
yQzss/d8xNqIVnePSZ0y3NWxIgvpR+ePoN2Spkzk4D3zq/p5ahezJBwhPohY053AYgPu1zJQpjOH
qJ8l99pr28EY9r1uovh9fjVxTn9xVDrtsoqo2pebTo6BHbABsi9VhYIie8GLA8pWHm8fCwKDvjOa
dI1+5ahky1SbwZkgD9+Nyi38OHq/nAKV6GW76MuUV+SwhxYyAVsMrskEZx0LhbT0qQDlsgGoqoo5
F5/lulKT4lbW24uE8sQvK2Q6DFJ9Un5OD+RPjZO18lyPmv9364KWlq8HqS4g0Fayl8COpSJvIFtu
hgaH37TBdQ8ixKp6bL+kxTf/acWGtZw8GtkxVw8yzhUqXj4C1qJuzbWeNBnNF3GLb5FeqLRbfd78
Up8yPedj4WxTWllsA/D/HChFOpkFVkcb3yfcVTyzPt6LVVeQqtf/9EwBkN5HptH59DI3JK6rEkIh
1HtL/gBPmsLtP3WI4rcHy+/xnBuELwG7o5d4+ljuX+634WWHaeiBLpNILhx1j/j7/ViJRHfxm/wJ
bEgrBBMNLKrnxo/XPb7dK0huz1/FwH5itDu9t21AqVwh/kbx1TV2MvTKyvubN16N1R8x4uwDJRHz
anATORZWq7qdDjd0haZUbeimBCW2X2NPhDmMGRDx6qJmlvvLMKTdrf/BaoB4dV1uQrRQutO5hRIp
pBG+7VQd3zfNMqXUqLIpnK0co+KQ8Q7YHmIE5zAUp7HeVFqC5ERlNjS2eZstjwaJdThLniKSH+Tq
tsIQDIS36tPveQi0uBHO/GdqvzvTRmyUbMFR/lq2tzou3bivBG/lfrEAzZGVby47anF6mGq6kMAa
Wd5x2+nQbM8gDX08s5SALb6JM/uaNlD9lbhdLk9OklZq9V2DAd5khro3xuFKPWG8pU8wz7Uy6Nlt
D4yyMLaE6JtrTGXBF4zF7SeDfAKH4qS/ouExKykZtdXT1nAQ3/4Hkv8JfzJigG+PSsuRI9jPgxP4
bNpLy5LSAlt2UlN+Bun4SzXLDfLeJvyZwVOMYD8nCSXiYSWW0DQ2yV8/P4CQ1ysxwyr90dtp9uAK
AVc3A81Gm4dMZBL7z9SmKjIu36V1GKN8usBbhOC8o2N5QvCctIZM2fM9dfbNEuESOrONCfpKgoUa
88eMa+0LyolkfQjoDJOUbv95Mf/e4B9Zmy7yDdaEVdws8nMDLbKsPC6gTubj4pfjjs2qy+KBBV9t
nk2dPztHwk0+43Eae8TwsMXBXiZSf3GPuPxtaji7onB2eSdjqWRR0cCI2yDsbR3e5LGdxRE/BuYS
PTZpIo7EAlkNBrSAAGMoOCyQczxIL9B+RiJd/Bfkkc3EEtJmq0+1Vq6MpO30KBvFWRExmg/CQnb9
qWcLhcXtbyr23Ucwis4Y+kwc9qOxOhltbus+3dN0PW99PQrUmUU4QlBovek1Vfw5W/t9HbyWB8Zj
bF3fVJhZ9eGIJzvmQ/+qIMp+1lFs7yrlhMDthC8/IKmN5ir1+OXth/cG4kptDuZyyMJVDI+WAiA8
11kOBNTCa+u/aVFHz4vWRrzGg869mgQKBkV8e/otBzrUEq6IL4bS0PcwanSnjnynqT7V5YIc789S
i8BIsAQdOzovLl/l15vzHsg2zmGZj8HxpVqgyt+YeuJtIN4r3dhuQFZYgoNIxiZfm8nhfpzHeW9B
2/LKeoZHPtsrAp/KZatYlGdINGNQ1HKahXMBNgIrJqfPLUJ3vwQeSMF/PBM7aLltnGpzDcU8lJSR
M0Rgm/jd7C9azDwBcD5vpMZJPCPi9NnE2iqia8elYNJ3SWYAKYdvjv+LkUn8kXHMALMQdwj3zndj
FucM3URzKmuD0rAHcnUWEdqHDx0EyDEcF3s0+hrMzr2LJkvtGUTLB6aEctekaV/4IhVlITyu/gqZ
YuRbge8mND6U5pxHgYvpe99eVMstYWT4jd02b3TK18GlFJVZe9b9/XZzxxfE2UJFSJ5l2DLsARMz
lc70O5wKM8yN0Jj5cUU43j9VjmXVqerPhpj8yi1+97dhxb1D/433q2lEczHqJTALMsMyaAjbzpaR
SfwOYu2iFO3BrCaBAV/MaXnxL9k5Yf5KTKeoC6ART1UmbBTKUXh9MpdKNYz5GNksvZKlvTQVikzg
IxxpoaxhREBWgI80jYKw1166vytsJgu7dyH6JsL8WUpKy167R/V/nROGASgCANPQ7iU0ku+FCXU/
9XhSvt6qhr7VOOELGK6XHlyYCQ0gi34myTKAbMklMNyphYJzo8VZYiChOyzftdflPDYJmVbGUYaY
7Ea5RdW7/d5Yl1fqsWn0gTVKjJr6cTRLBlnABm5QBxDbYnVxz1OKHVtB5CAzvhJ6cSZo/Tz8YMHI
WngKsxCI8PSbkagWYRh0RH/MzC0OnkWEd08088sA8XNfhmYTxQuDW41zeZBopeTacFptKM4B7OXO
23/ia9juI4vKg0zTkjltKf0qkDiLIqBUAiui1lBQ8asjKNPUMfI7ENgEkph8dtE+ln3pW1uH1wVz
6HnXmSn4zmDp2yVZOSMYCUthCjXxeMVjwsd+ofyUhIE+3k5EHQYYO4zsryA5PCgnVGaPUMt0uJyx
fisQI0sFI53lnSdCwZ85YhAwcoQjCkZt46afNrp62+SMG0Vj4awgFAqkPjzdTIjGjNS48k8t4M9e
gQsTc0+bOg831/CHgItSMRk97L7XAUs3p3z+jVlyn9iNB3hQtF0a/nZ/0HC10YvAKPtKsnnN16Uz
b8K/QqdLpCYs/1dE9BwMw9soQxG+pMBdxwsJnMHo+AN6afE1E3V8h/8pTxKby1GOVXqf13k2IcQC
dao3QYJcSaKzfECW6HSfgLy9tUX5mz2FdZNznn4QTqHB9U0eAYGAmfnJ/tlbA8PoiI+JshFDLODu
kOyJctlPFrmhIALvW4UFyMoiDbWsdqq2KY9EKq4wzrZf1oPuDDF+erjPTTlFU4jB1Jhr7SQb++Rt
b5lYlLafrqDUmBTmzmajR4FvO5abak6ISZJ0E/NpgIGKpuSfwgoCuTmc3hIAm0T4n7BUED/0iV4G
E4F9CUbWd0/1ZbgIxh2WyU/e4mXpDbCeyttkkM/6DoukLABborkLW9g6YG1T9Bwn+XzxVlICDDuV
+K8UFA2+7evoA9v857KnS8nzwDIyqyB9T0uM1n5F1ACDFSnC/cNJmih6VX+VntBCamCc1I9Oy0/X
/kPmRKz+CLY05Tv8jsYz+IZKliIn4gVsrQYipwt1aV/TR2cF5q9bdORa+wsi1oG+6Bni/qWqbNMo
IcH9HxBYwdXY35vVJBiYrdcQ71LRLKRDbhuL62F8yHD+6Eo/pI1MVXLIf5bbpPgceMdWYBlw9Uki
z/WlS+v8/N+RWkisAgxcY6+1P60y1GCwnqi/NlDhUaVXdzHXGHsO6P1p6MevPLJbFN7tjlLYevmu
3YkR8lk9BspSeh+LqW27Ed2NzmBpazQ+N0oEwly/x63OmwnyfLXSv4sH5+yW3dSS2VaY4T/0enwy
C0/AEFC0Skw34w1Zi+qHEUZM5/fSADkTMlEKpVFcEcf1kMtbUuZkZbbsyVPCF2ioqQ7+pnNZcRAB
xseTeyf617OYeKXjPB/KUY/+jxZNkcbOT0Dqvwp9yxCK9iGnqXovz15MVrMyekKB0imJiGflDAZs
sHjYtP5hBnOgSDL16acxw/ArJAyKfFSw/kJNQ44tFR5Vc7Sw8Eta1+SHVw9l2iROcCgFR92B5n3z
ts8+xvHVDKGlVxWMlay7J70jE34iuOzfyps0Y68kKaSpEeUcAqXHajr9NlBq5iplRFDGmxqoZFYS
vyGtNPM7fNZF6sExDyabN27hwaWTSe+h1vVasla7NR0JwYr5mCRis9+IMHxMv3rfSaH+oz+JuT8N
fyFe+Bp4joL5Ja0Wd7rdC7I3CD6g3hQGx452jjEXx4Uv1AB8qqpLF8c1Y2qWQt7hpeKXEOchhpGO
S+orRwlpQcyw1CLeJ+QFrBpZeDHL+E/6+v6ywNNYcHibzrmgl2s7u5jKIeECBRM4VFz0Hn4B/ByL
e3KfTQ3qu5pnPe6hbMFgPP+rEndiHcF+61syo2XrYtoy1j9afxQ3rviInywDNGSDB4fURiAKWh+N
2Nhlm7xr7TyexJwRreZrj3/MDsK/VJDDYNWA6eRBqr43ys2QxuLeHD7At7QmMeBO230EqyjV+jMt
QEKYVAQ+sDkF1MCM1ijHBxYcMaB53/Lubv5Y0XOJtAAUkccdqNApKeoPZdNCMkwuuiZ7mjxXBqiI
FNA3314Cp6TFLFJo8IavyGPi2p9kEVsRBQNpNpt/NxtXGBfsWoI+ZU1YIIxkqZiSOqkTYNUAeUXR
82UIiubmn+cddYMZvfb8V+2jEBrkTXuFz9133EgfyKGuA3yx4oCjB613oPwoAlGp90+lHBEIQhzx
aiu3L32Up9Z0udXEGjK0j01re+68KjTTyWIEuS3aC3RcbcuixqFGXzAJ1h6e9ycq7qz8CiC1p2zb
vH0j3QUG0fvmWoKGxBaVj/HmHYjL4sHOJAZ5zM6n5mqumW2WA4+OVzqakLQPnqSPRwhq/eYa1CCo
NIq/eiof20uuvINLm6LF5Byy5Xl4Zkfl16yZLCfWMoN6iw7O8RGiNv4m0g1fNYkgtppBoMnKSQFh
GAa+U141djKlz1PPQw8zhAzgNcIVqWBCX3qVxa+PabBRcd5jQvdXtRGg6QIMSR4FV4mLDKucSbKv
SPLAL5EKiqbrEZCHwWRw+4V2j1dwV+ksE4bhj+XKPBsRW07eOT5CzFEWYtn2zXfY/ievJoiuWhFf
WHPRJStBGivhTdsK3Ed8jXAJHJ2UBD/QdRRyKZhxOttaOMSL9SW+4AVt1FvWz0ONV8p5rTQZg5NF
aKlTHKA5mXq9XR5CU4BJfMLbJWMZ3NALBXseOxhmJr2d6I7t5m+teJh8RUy5QGRBQChjA0IIKL+D
IuDecg7YbDiJ5VKqlRBpoR2gWAiJgRBVGWPo17GVT0dIMsGnQdHOqsooOdp2L9F16vplX5qkVpiX
IzDH3gBaO1k/tldlPUntIfTdV71KbwT3W+TxL2AiAfz1erlzD050S8Mw7RO3mBeJcDsblY25ddzf
NmjERzmdD6J65f/FW7BJj6V5WWN95fuWfr4B50Mg7i1110ROTx2MEGrBaX6/t1oIicvh8JEqo/aU
TCBF8bWbKsWhzZw4LXIemy7wFTHPzLm+S7e+eVAnHCRhnZ9+YDMJ8PwcYv95E9NfNp1V2wejJ0jD
iiHLXOq3+yu3abzJDiZOnVsHxnyYfvfs2NjLsE3O8P6M24mRKBAY+uT/Zu8SchEbG2Mvk4GypUBn
zD0C+2waBACmP+By4B90tIXCljXA2BR0gLjzjojsRW58njs+1AkGc/9DVy3JpH+rccVCJTzJaAfu
mHpky9PtW2zeshLXdsz5tYDZdEwkwlh2q0TWvPuuBZypQoGYxA7yQY/3+SvwCa9XIQFHwrqsK3fr
uPiawy5BAC8rL0EtxLuuujW8zz1/CRCIi70rYbhSgR5Qo2usqzVyvfGT0KD6Yko+mMQcz+zN+Jz0
uL2tJVKbbD6Ii3dHNhVFMIJgvlMJGLuO4lPLR/Ft1ruIwzCsNB511uQfPHhQujo655o2ShSFbEDC
2ROYK699RLYMOX7MsivI6PTeUk5hWbz7RlUjltAsfV+C4Z0YlBgQ0igiIt1JoTAynew/fPo1ITGZ
uAZy5QK4eLytANerx/4kz0qn4tLanrKnWcE2x+qAvRQEI1L9NGdB3jo2VCYd3CbEDO23yMaYFvbu
6SLDhC65aGWbYkUfjjtP8UWzcM8Eq/5oFYwffpoew9jxEX4/DSw1cA5ZAGbeY6sq2R9/DgwpATtN
Bg4cUpPBDBy+OhJ4JGCZCulG8zNcwTTLu+ppvAtZ2QcY79k1iHJtuDhBsAGjOfW/V57dVBM40UiT
d+SsdmvyHdsONm4IJJPSZ3e58wfGogkUfIqlw6BHgHqA876ThF5gF0UPlXL74lniVI9NIR2wC56h
/l4T9eybPecWmgtgFlJfsbBTbSp0HzPL5KDxAi7gBhEqunDfQK1Gy1JfKbzVcPB+NSamAe1jW7KX
OR/Q6bKAhRs9uPoAGCbbSD67+k4YpIna3ju56XTadTqvluko8ema4krroLoA1NJEleIhT86Vrz2U
9HDnfJEqNszlGlJW3vsRSurEwYCGvavTxRHoq96Q6CnLMDKMSHqRj0e/XwbYTRxEpD5Nzfyj9vEV
Vq7jRf1Bpg0UchBc1rmMHwRCvJMDJDk3JAnrjBM2eD/lbqEvESqPg1aWn84bAsUwwDszP7S0bhwY
pLWu4gdLXoVlVYAzPGg/ThD0KN7pVoVUqZl+dJGprw8og8EXRC/v5o25Qk6rrr4q68XV9boXi0Qs
iJaKDIWMr0+2Un2tFxlbN0FDDT0DzKWWToXG8NC/zqRlro+Cp80ujk3WFo8QXXGAVYz4BUxMXaP/
28FtQbBGELN4WRqXs5pk2UEw82157ER7pexgwqobtyuA9p7DQ2Q1SlNLMmg+ewjMQmM+9zB7d413
LRYvs7HiUzcZtCwjkX124rY9YBGbsG+yTRCdQlihPX5M6uKIx2XnKbO5zSX2cTT8BfvkiKSG8cKt
M7EWO5Hul4MehSrKe3x+8SpPCbXIOe2CcE4p9dQWgDS92ogQxZUeRFe7oUtJJIcYpAm6Xf2295HC
NrHXpgV+dB7CuBi5KcrdvmR3mHw3XBFN5MztVdFS55ZvWoVbbydpNkaqm8Y8UL9007shIWXyZDds
WTKn/gqnZdA27z1Q6D0DJGxX3pOzSktQLz2lwMFqfFU9Q20OgN4PQXVYxNf4NVQ5ZnL3lK0J6DkN
VOPwgDudemKKQEEw8+UcMK5PNPVkSrIzklmfATwTdvmhVvnkG+q+rtTY/GvtYsb9wr4pmwlrE/C+
+KnOs9ABpkN44yS2xzJX8OjInxxBHe7+xdutE2JwTQ1HfrAsm6ZF8V1Hqv1+tIOnixlgD46MbVzK
M9AqyiTIssw5QMx691uF6EbQv/62mM53BRp9q7Hk4vo4iRSCJmRFhW8Hg9c4gRB5lEM5gKPDAifI
P05DwRFdE9yBWZ3SPyP7AVYvFP/hw5o3eIX0ivcPVT56gOQ8b2PZnoef7fzobwTnzJ9735o54tIh
I4PnbY5ghYkLAEVvXHoJnn77kouy6OxPSc+4mD56XeGB7SvXoj5AfeijUM0dHKO0w1nZ3V1hcE8y
+Vps6Ss9E8UIv4forN5X5pMdzW9i9pR/9j706DVdSCl/YTmi06Df5lpXeYj2lHyK2aC2wBZbdYno
yoeU6j+gzEjEACj+FFgRIUY84tarWLOm43423A2JPS/xfu6yMnpDVdMK/MIQBWaFzbBf7tVNRHzV
ZswVBqzbFU+G/F1rkhGt1uqW2nEh3REpPAXFUT89fhfWCt9dLYAvtJpFmXiLZLvLL0gSsSKMq+ZA
M6U/sGT1/J+JH8moD72aeRjI76QA0vgjJGZUXAXVHpWsYjEYS3S1+fLgMZRo05GddGaXXncNvYnE
s+cRJFmM+pM4L+aTxgwxSPLZPypevJofvVpl531Rryc4mxUIHI/Pb0g23/Ve/OMPVT4k4fZ3tkfA
8WEkuH27gqIFbBGMmEWMxJaSbrHXFXbc3adH6TBNw6nP9hrz8aa+o0dTgQJi7l+wj4qgBsqWDqUy
nmk22upUuJRaXw32idLwExzxrP+/zg1yABOW9lkz3M6FrFQz+hxTRQ1OR3cO/mmylBTUeXZ9vZYc
1haxF9Ije+UoqkZBQTxbeNZWu4VbPR3n8+6Rz7OqXcSdCDk4981zoXtr3S1hTCFBTATQBzwRtilE
OUZnfemJfcL87KMYQqmBeuZa8907ustMMsvKt+RFQ+qpiVSrszpPMeVjvK4ZzT2b/VpY5U3gfb73
STrkCPLf3lbDC4LmprY77OuX0x71OZS0TsGGr/ls1LrvnSUQzaEGfOQQEL1GBXuHYSvsX5UZE5aw
u1XKmfCWViTi43l8Y1tg32jOiZ6PfS5K4ZiFT15XZzrzk/Tqaaqqs7vDKa45TM3Pou33jjpjF7op
Tj7PuFy6FECc2miR84bhitbPrqiGMR2+M+4Cn/yugLZ00VOwZm7wqVmos7sB8t490yvb55L2g+RD
XFpvuSo1DOVWrG8YP6Yc4bs5OHBtN7wZOXSWsNoOW2LtpRHvcOrZYzd7lHNClSgtqo/zlGnXcu9q
K/9KYmyq9UmhwgtE1aZecbagc/Qu3J4vjqsGxWVkamQqrWhQsDeFpfsXhmN6nJ4jNTa7MQLfnIv0
5rdsh6REuqPZoFrYYLV80Fm5cyjyRwaVmNJauLFtAPryXdEr/FjlAXd5ZVSQeG7NH6CVkEI9ymTC
9paKxsK/QCbiibT1HyCwWKJm9XauVMfVneb0SNWOumYLFLcjEKU+zN7++ZsW3GJS69p3AEW4EX2i
zed1sHc6q7gsiwE7mQdSiSfo+KNY9UoVRHNTxGSLSR/7Zy99VNRxbBDKFoxgQfFpoi7SgnIaXT5x
DftNRm165K7W+IahMxeHfIeJnwEXWE9w5Oj1aFhmcc9rLvRO5zP4XE0K11fSVbzVwhwVbCy/kvrF
cemIqHiM9D5XcmZVaMfayO0Y/1mv/0gLy1KLPaOZGNOQK8Ks4ptiik+Ne41boaCbqjo2OYaFo0jn
RtvZcmLkRhB6sH01NTnUziouGvM1PIKeL8SHvWcp+o/7Dshc0REljnixhczflb8cH3NlFS/0ZCqf
9E1Twy8Z3gllnvxumosYtyaFc0qqrjQA7Vl2eH4F7Au+vI9MkVNy5DzOf4gwywEnBqS7j9ZXDDfJ
5iAdLqKt3K00zZaaQoigb60O7RJwXtPkovKmDmsQNqqI+LndSq3f8yaBCjOnigQ/WO3+P4u5wWRP
AD2J6GODCLzftaChtKsegxZWsHdzrnuv0wTiC0yAMqU8AphsGzBjCbGAd0nTPwXxrgaj5Zyrzm23
rSQjZpLJmJH2Jx0v/r17ehXwSLZFB6jbV7TxA7V/IMqY/1VHTWGQJuQdJcoanDgh4hflVvGhY/4y
VxEuWmH4TJwGkwibb+W9VNYCMtDVLGYMEdmjVun0qwASLxnEaGWHEGgvEVkl/7IoEvoaaZ1EaBBi
7qiqzyGuNw3twznxLpa3jGuXuMxvP+rPb+v59fZilAUKw5EfNNnss3oBeNNhxGDpS4wyzJoD/Un/
wX+x0otlEgmjBs3grcdynIN70eFzU3WmZtwZOiqvBq8soqZNIUfq10mxYS+4lEIwChvASK+PXH2o
4/WVms75JlTn751WKGjvHxKenq9IUHJ+xPhNDBBZgzhyG4gM4MRQH1pZ5my2TruIA7sVImMaEnmc
eezHvxCikgUR2Qu94utaUcAOMzle2xD8oNLkqxWKS2F+i3uDtqhkkcayoRLlcoBE5vpDZkUW9sat
PtEzIdDICRnEKdLvNN5OVZU7Yhl/9m6AJaerU+JAED+uIYazebSS+yb2pn9WTJB81UJE/Hz/3uZV
kVVQj729dULaJWi8yVq/YhTjgi16c9tt7la+WxuTxRC3W7WKJnBpk+Tk0Wo29cSxE91vWdjppYGn
gbrEv63vkwso2qpKpCRQ2RQd6TmpZTduhS+/m7kr4ELdLsSCFXyWrNoy7rl9PproUd0xZxKV80az
qcmSqo70bNl2KE4gV0xYofNSJGU95iCB8rIkPqN7bDYJyx9qvfKn5PiBFhKbOvvjThP2LOVeGn69
cKtUxW8xW01rCcaCaKdhH68DKOEYD2aJGEOp/taMyLSS9aLNYHIYb9rSmqlWW0P6uvnvWUNc3/pj
0AoxqUz5w2gMpw9Ef6y5V6YFMaYD1e93g65vTVmJFoy8cR9xuYKVJCsZeJIPXfKXKwJ0Qk0n8+pt
8tQoFES3ZRS/M51o9iC/XXh05L6aSYi+q9IOC1+L/hiMNSjpivg8nP355wGvGZfGaLBYPXz57gXg
9oMKj6KXzIngnqoxIBjEDOQeEfIJH+T7pOQYRhseQW6p0eMWx/m1SUuoycbQscRVmDksOlpGvRzR
XP9qNrpHua0EacLcrNVu8YrS/IRHDgORs8D7uejNWmf16QoKGZ7+mhifjXknPjxxHvESL2bS8FdB
HflhCPIPCejE9kZF/wmkt2aVkibmINz2w+9HPoWVK19w97SHEZIvNFFe3o+Y0eNpVtulwoTKrWYv
hkdLDst6ejADBVY0J0/wCQpPYngz3Ttz5/Lbmf+ojjyFSYClGHEdzaclYtSqT4n2QDlqIZf0QiZC
/z3JVSCcZpH+7Qn4d4btt8KoLgJAT4qyWSwlTPfJu06KNUQroH5pTP6alUGMwjrfCFa8nOvBQGLC
9dvoSiKfMrbK/2SEquuXb6ZG7Tp1wVdKJWLGS3kKzvzlRhVzRwhoOWnbHPr+LA0/FDcUnwZQQuv6
z2CXI5Y2+OCWt9DHeWVQMGjPguMMwRQIyRNI83Befd66thL/DHHDXcKmfN0QCU2O1NN7RD7ZJewi
FOWzytjYWdOhrWh0DugdeWauqcPmpLY2bV+GwJKjhqtFArMNTSX7n73oYUc76Sbq7A5UBk3fIp7o
1LftzeLIFpMB1nhhXc2jEuIr7G6SJjQC3kNxYcI/iTF4X6X3JcnOcbDJPqaw2G4a//zzYaC9UOgj
phvQ32zeh6AnPN1GWoIcqfA1ETXJmpbSBEHkVAvuskFbYrqHQ/nyoFzi0UkmW7NURA5wfesS3X1p
5bwQfefRSYQTwLhzvi9TsUWQcFdT4BZTNfwdud6+lzxa8p+73suin72jsReI3eTJJ2nfAkoX1MYc
fRwR4TTRO3wUc53+EK4bnpEvULKRJQk8FghnDRqx8r3b7YRv/qJJlQmv/yfLjF4VqLFdznAeX6Km
ClphTQrns8kQLS7oUrHu1Wv1NN5iek34aKpbN79PDGwjnAfAXawDTN/NkFd35pSaBRberrC3Eok4
JNncSh4JfrUdWj1n74XPms3rPlOG5mOSqtzOvI+5SafS8ntkWGT8AvN8/mRDUUqkzPQ/+XmvKRc7
erxRGRzBlQOI9j3eTfvWGHiwd4DDegWVny/6UYM6Rb4pmFK7xHkygEoFMchJEVrH1/9kO7H+O/Ou
ZhIi7g3GrbyWfpWv9FbLwR70SZG2PYoW+YmhiolJEYp2HiAmLJ7LcB27s6tBhUE41huQm3eDRmz8
xiUFB8Qvbo3PJKoIDYo2/oyD8KN+qxvHDeqQQA5lqB7JwmyAc/BAUv6de6O2s+o2/qVrim1AQayh
TM/4/JTXoODgsMu/bAEfGqrWDPd0itMdkCeiMrGi5E9puIeFs3s7+opnjf3V3LOdKLckxUBZLav3
onCcLW3uhqGU8pyh3ZNZfIcKveSsaxTwLuU7xLlU35+kXoVJg4iCadhcFjulmZgU28p+mWZHe2iB
2yCX9OSEzh7iW3/n4TTPPk6yqqf4o9ZTgHo0uVcg5VbKYDk48XIqKU4xE2ggWfRV3h7ZKmsZsteZ
7CbVD7Si6HFe1x346yyQhVE2t00bAwxwBnhyRg9BSN2J4G6TB2bUO+8bEQc27vVhdJU+xrc8n7ZW
MV34I/qALwJn9wiLquUf67G3w30dHL1EloI74zXkQhAX0XA5qDa46HAJ724+pTsZBwzQzPyYiAVn
Ol00YaPE5bV9L+q+6NVupYqbTeR+Av/I9zQY/iP0zieJ+NyQwjb19JT7Gi87K1lKJudu7oBADQUo
e3wAmWeZsggo15P6I9Bi4g5rcjLlFJvfTSP9MHCpXWnK7w+sPzTrZOxgntKrQ9MyuKd88/IlRXiA
3zBBVxpKdKqHPDdbJ6kj3xkblW1xMLgIKtdbEMgROE47vSXGTqBF5Msq6WMIwGqMAn4sYBZd08wD
H9+MKWjVr6FqoQxmfVXDBNhOk+4GEtyuSAKlXk8Z2OgHKktHLD+xRJYDuesETvSDn2UQUnG2nCxs
GYv3gO1CPFVLtcB13J8dcxur7S6VOSDta5SJoxLJPqXYBmDi5kouK6D1/QsmA8rS43vGs0zj2S3C
CaQ2W2nArW+W+upZv1MDod0D1rlNaG0JtjM8Yx30fVVuFZaqMq5ifSOFh1+hr6+FqaL6Hbo5YVad
t2ZaXI3ThJ94VsN0koVL8z45wNdXPoIDs1mRT81Tjppet417dAvkljhYupWTO3kffb7/1j69btOF
wOezwBlx6XmyKtvcM1jcb50pWO3OvPWncK2D6+xA4rNgeOVI+J/yF2vWBcsGkk1h/7+z77/wBpVu
+nDgdH3JpX+0GIRpQbXlHA/gjBue2GJHttF5+MBy0XaiK34zhe6DU+aMQdOxI7rUps7IReCyNopm
ITw3JzMUYKn1+++h9kOxR2yTHbuIS95fkh8Nr0+T1hXPuP/LdL9QXh9vzCLj9Fy3tAF4Umb9hAoM
e+8RYUyEVav40DN+t6+vuhDtK1M6YJEMDbKjwWi+K0r9K1ZQngUlrrsJsNK4QWiTCqI4COEy/WG2
gEZ5lqD4/kO8q0EtM7b0KwEUR0mKFSsZYehTUnNL+KLD9APul5OGcY/8EsEjKzUkIGufU694Q+mp
6GFVZCDL50C9k70gd/JcXMl2fL+ELefUoIMwqg9VkME5e4Exq9WnA+rI2Ed3+zi7zJYPrPBrCWP8
8pYyumpxDAFI8R6MUlng1VSx/o2yWR9m+weSGgX2McADuyvXHjghwCsOfjAfBTjnLzIZmn55FEcu
ybUgGFofbazh4XqEFqAKYu7n3eqeU+ro2KnbMD/Mc7P3Jo4DPo+xBjrkRMH9XdmQJZmz5ePynpoa
tJT+Cf6MJKPJARVZex6HV4eyB9lTrGDo0gu45XxfHjGGx70elWcY0+/QjiQRQltzUgvKilbCvX9V
bnmAudHKnFFgw8szldvlZinwgIjZ6zkigUmzq8c4rhkeXajSMEueVoUlgxUpMm9uH4XNVJGFqsw+
U9U/DFSoHIhn/3H24OVR15X19Zr8ZZz16InnOVFq2zXUrpAoj4o+jVFtxz4s9iw7YwWDVJxRyXHu
csYFScXHFTd4fIcccFshWW8AzvcjJno0FHCmG115qDhmkGe7IxpcCncQx11Tg0sfqG4lqUZpBp9e
TRARpNcyvGUDvQgEs3vYhDmDhY4t1FDN/YOfed7e1xX1CNdoVbkCOMaCSIk3WH8+fHljx8nS2U4K
MU6SfRFU27lnb2PRgrUH58InkokImcXFnOazUniO4/f/6Lc8UJ45q6IgO0vWItcvGhcVEEiB/XNP
oAXjOuHUJTODrd98g9wmq6nXR4Dee+04FsdFbUYJDX+wrSSpJXf+iQMXZjiC5f+fsf744Kf53PnE
E5hTsnsJ1o8kholmyo846XTGcT9qHwnku3wlU9UGiPL46Xay0R4N3LnD1FFs6no6Bbrty38Wqg+A
GvSNtk+uQnAKDhSwRl4uTZ5PAjIcPZEhj29CY00pTbeTjyYYJTDqMNiStDYGoFoI1vaPLQ3XazoR
1IEs3J7zsd1VadRNzavEeisITepxmXCVValFF0EUwbZXYVOVRuHEr9wnL225YO1KTDJL8vZRu2t2
IHRz/LYsZhhPQ1WJSCaVj9oPZabJjFAIbn4ZSp4AUwG4MNch9tzZVfLAZIMYRO69qJ7EotLsMkeX
AdnCmqS0YTBc1KltCoxmZQPuVmpnwNVFILpxSgpGBL6ByzW38U/T71OeFe/FW0YrKSd7QL5zzYOC
LgWagujBVyY6b93VJ8ZDulfENUS9JqhQ9y09QN7THAZAO1vWf/Bdasskws1DuV0SePiNgHKU32yx
9e/aFkmJooHr8MVwUpAaGyqSeoI3rMFk6ixEqs95Tns0mZKApO/UjO7FZnf3BIuY3xVjxXd9XzQd
2NIFOWIfPC3kOEpWiBK615hoTNlnZ8pUoyN8pe/QJuH37kspezrHAsSo3EdbWKAja6knvgYcW0zk
x/bS3xif9ZCgEcrut79Gxa+HhPENGBGyHa0aaHYUlWylv5j72SIrrM5d2NoAX/eQzqOaiHkVCoKh
OKayZJ/GokQYEahcR5SUNX2/6T0pELJrAAJAgeSuyheAWfgzud1pORo+AsHCECjSJdro3E1xdTcV
Rw4aYP4VGxYFtwK1pW8nN8uPSCfq9lUN6smzesx/rdYUTlUWqEJB+Oxq6vnWtQSPlyTRsBBs2CtH
7J2muGewQmXVapFS7+aJmxzZgwAXoaoug+x6Ej9K3gkNpH6G2y9A15UVRGEcH/MfppfY4bjSK92S
5J0HRtrndmm8XIKjnWgzGa2YT67V6gPjBIo4vhyYNvGGLqug6u4rWoL6aTyjDE0ocVT2K7smudQT
hU3bXHDDnFpT2m7TyXmbRK/QZ2GYixTKbTtOyU2LKco+AQoa6ZKz/w0ktAjrwfnWXq/ATM0m4dg/
sUyrita2GcRGXygpWKELTeWbR2/CxD6rnJVXfjD5dKUk9R3dYNxEBs46VmI3PwfyLSo6Y/j7TCjQ
KPfc4Dg9+hZ8oV+FwUJRBL0ruwnP98ibjeAMdJq8ZQp/52y+KDtUloSAPR1KQfhFO7NPz9SWfD15
G4ov5nw+9LfkYUG276KX2Em8r0jfQ9JT18nMxw9fXeEFp/0kL8c/FQmkcz1CM9VcsoFLuFoAe5pp
O8iRSHBU1pClS8Hnp+vUDFU0fJPoK/qC/KV7zXp+3zzeOyw2BNa+Bd+W8QYstYnJzYExSOt3niPz
tPPm75QjzfsWSs7ENAIDF5+P+kXTUgZt+NRm7g55qgb6A+hXHtjZ7Jvk/+jq0nmUo5fMWJ+XCIJf
TQyKC1YaSehevouccDW6kwRO2Wx2PPV3MFRyRisNzTqDmCkMBNFqX/r1XIZ3vwBIfDtbT4hj3vQC
95140L0/oPluKjWRecV5NUmUQlZxpA0N2rHtQD7jl9Dva0wNGTswTxM69VoRHu9U0AjZ+NHKASfY
sTLQI6LAYhV31kUvwDqK3JOUU5PVmsYDkPPEcxhadV6OWNhpmrSPWejEQMpP9XIHag+ySVHOx60k
hzQMD3Qevsf//6dRM0aj7W6DKBCeR4kBXJR8+B4BiuVQtE4mFOjnDw+hGvsoSuLjbeM/E5ZEZYrK
cd4N+BlPY8ru6AXtn/2waMq0ATd9e2VH6HY/nv8DguSOlYEOSrQeGuaXX9Y71bJOrsQj+tnv3TWB
juK7JF3sI4ClJTimf9Gmf7j6wXZ6TpQ9qBD7seNbuB5hLw8HGd8qrQiqpAXl2+RnLVaSWG2VCCIz
CEx5/DFvrS77rZr3nP99PWi75Xo9dYWSdwzm7yrVmI9F6RZ2hFMAvvtm4pvACMMS5YXloegkniQK
XF0IHLQLI6NBONj80W9iCZRPiTX3MrT9KFhnClLXhtZJk2DPJdQiYI24O2L1y27CR0aEblKcJlT9
CNc+3wno/Tw6Mrh57YfplRVM2w8VftBgFcH67S9qqpTmAeDTzzmeNqDiI++bZTmBUn7TRBiY0oGz
mFsIireMnGeJEiGOMTlS2BbPCLg5P4W4qXjA8kb11Jk5UpV7Gg0Ph9TqXf5/RcOxDodq8BiYpFVI
UBYHYJal1zdLxxF/8PDtoVZ4ODrkGaRSioCvAi2SKfcy4cm28nct5Nx40F850Hpn1III12c/HyDb
wg2wYrvi13zVNy0GY9t62tKDlz00FPd+fuH5wU2O1zcqq2UWA2G/o5ttgDjn1P5Co43N4ZiW/6/r
GcdzvpLlGI9h51rb30R2XHVia17EfmUkROXcs5bFP64zr0WE1oAgDvhlkhrmxL3SO9sp3uyOypPv
whxmX1ocy+w+S9rzpoW8GA3o8OspwUItjoHU0SjCbluz0gV7j/Sj5vIVF+desC6W6w/BaZj1IweO
OBg6ARZS7XO7mLPoqOt+mJ5/c8HBJz5o4kZWLNuB8z4/QQPGpmoqKCMpN1RFDtUvly8cT82Frn7D
HcWrBIUNaL4DL/BPbHlMA5C4YiqTXafyzvhQ8tiqutumzfRUOjLGNtYOu1Y372UlFEX0xDFxcpZL
GAEWgR+jjf8IjZlOE0g41h/zeDswCHN9ez6d4DSgmhdQ7spuCSgBQzLHt41+0IzQ0bDzjLypGlCT
O9jTea75GxsQ5wO1ihumpf7i0I0NP6gAsa/xi0gQxDj2MMwQcNfYgNBqrvYvBCbBmdMFijsE3DR3
4uwAfnZid4QroTTHCDwBKcle7pOqmbppl/DtANUptFtsrjQWAkVp5yVPsEJhWXetmu/asphjqxRz
8/DL23b9+7V576JDqwtPOi0O2Jqjb6eSDOg5BTxlYIGN7wfRxQdv9TlizmkRSGtFXJeryR1i+Gbd
LyuZgqIdyt3l3GOOfHlxSOlWWJH/W/z/DmXC2sgnGLUGNvFgb7I3rxSvYGiFcp5qo9b30CEoZO5r
TZ5R/JidTjrW+qsHIJqqoywZwflFG/3U7cevA7XJhrkb482CNUqqFpFlUzSbb+BqsBGiBANlmtf9
Pk4i0XiKUTrfls6vxh3JtLYQgLSH/pT51uSlsybms01+8Oa2CmEGgrAFM/ZZpJEFGWDGBwFyOoVY
A3VUq2stRAVpwa53E5gn3F65JTzZG+b72HwXozvJ80OXBD/fUoy4mrQcuuOuLlopQ/Hv0RPG44Zb
/Bud4/ChZmik2BfhQYVwDRjGWPIWyw3UTkWxYMQ5bG/oTaNh5ezFAXQDzBfBxvZKZarw3Eu08m83
2BivIHmYYAlMgqJOjWoybg7VD4kElGYkJjVTeB9hU5EXq3C2giAoWpzLE67gl9q6cFy5fbe60KdA
dMbssNUyFqPSjX+LkslEX5TaY2Cdj8mKMC8VhIEp63b+ugO7XWDvMcs46Jk4sJwRhfbkKZU7bKTG
iK8exSgjt8M+EQQH8mLuO+zfTBaYMsd0tmzs4TFWVXyYXHbrYGUsdugYaiXM/sArJtn7nj2T6WNy
kTqQUe7gqMZEhPytmTGop/YifcpTtZOtca3sQtGfVuaeZinnx3jKGnWIMaWES3ZqFOtQ+NmzpwFO
sKFYSgGY57P0jgv1S7ojtdaqCx7GAJTAuFhKs+gZ53KQSCLl9n+DYFqrk/57MN+GlmrI65WE/7Vj
chn+sOjLXBg19PIkdnh57f5iSr3BgwKOaQI4BnyWnOawAal2NDctRsR/xRkxxGlt+/gSGf1GoqJM
oUynSmT3iRFEvPUVONL60gcLSeH/gd4CtqncWhDgB6NTyM4w/n4qczo6u+7DTMzD4QOELz9v6BXR
81XporwUoKbcNVyRgqYtAM8wLOb6KvnXspzYQP6wRcoJmsSdBRJdFnHJvtVXDNzHA0b/DaU7orGF
0Y79KTPKPbSbTM5C0Tx4Izs6u6/Xi7vZ0vq/H9LxFYGrXNTWatJBrNBMkw9cypDJvLU58Kx6dYsd
y/gR35aa87mgbMh5GM8ils7zjv1mhcIF8HNSZOpDWy/9b891DiXEYDdYPFCzi+wgMGbkd1+L3TcX
In93oe2O/KKLv8UAnKS1BB6ptZWm+r16ZNDrO6UXDdm5XnR8qvaIE53R1ms2UFg6H3xtZ/7SrOw5
1/JAkXmP6lbiLgyQw6xgA9/EvapUisnl3XYInEIJbTSJNlZLn58r4sD0jmQqIepkQEkjq+ZUKLkE
Q0L1QPvxO4JA9jxjnL+9/XDCQ6h7MfOet9ohPPffgDfi/uJbWrpUXcDXdiSsU1nVqzOqrJ6VfEMH
sfBc5wKWraxkzWJnj6DOOnOvm4LiWSvWjmi8JeMR6G9eMmVPEQxqM6LshKo90iOJwflaLTqVpirc
2EPevzuMVPO18AMBXGL4UPX89xLgvbzT8Kx4popKDJPBfU/LIf8A3xIvqDUPa0J2Q8GoaUneFsvc
cYhSkXFP4pUb5K24qXUnIF5V0fk8R9pBam+/a11eHw3RbDrU/gPZXQZgMDFw/t9zHrtBJQ/qGZfX
XEatRRb/celyLk0nuav8yIeL6RdblG0VifuhwwDvMuLUVlw2EV9rMJ2jz0nxGc+nxPZX8LFHrpy8
5j0bfjguwCykNbsg9QYVR/NuJ3hhqqxGibw3MK2+JzY26TKLQgv4VPETC7RIWivrLlJEpRZ2IMQT
62OjEIS+5NW5S+E+hpVPInXKy9YhrZFlBhmadJnG4fzREboTqWtdOp/QA0kcONTxuQZ1utQJcp/S
qxIg1TNlhYwYV6873fb4d9AV7XWT35HHc2z8wa7YAePuSY7m2ilaeXfjSxcbjlnVfgsXnhWfUkop
+NtJOaUjm8ECyRjc6aGbB3qvDCkrNEKXQVC7px86PG2/Za5Y+swLxtb/mDecEjGqB98f/Iu+BUWE
Xud5L68IZF9WGTmwDsIzZIUfr73oQmD6n/rPI/krLdECOdX6jMPTB7U6Wrmaw3koRRp/1fPDprBA
gjAkN4J0BpvwG2C2DpFmebrRjW+QoiR7LrbNOlJ9nnm/s1upkWIMwnaR818zWvq6YvaDxN91KhKG
OEJ40sGeNPS58hxTjJ6BwVPYouFfCi4yhslL76m2LoBvTlc/f4yRaUzV8pZS7Wz4yMmsJBHP80yk
jUtEV0DDqDhRxWhBqONlHYhkGhQTeiqNBIU1p8C2fKE/6v201KMOrmQfVGomysFbyC686NMLUoUD
hGpbvMqbocp5/7UzdPzel/25utiw1E5xRj/EFk83xSbr/fliKj0aouUVZmzgKKeF/ClIsyw2H0WE
gdhEN0vfNp+6TBRk5Q7dxSxclSGdCo1OnPpxQdwvfUiHdct/CR//T6Yor/9w2D95dXI8Ouc1bNCU
nz8nMEZrtgzUx8LSKk1BEhhO7o/KYKa2+jiiOLLilt2d4vowB+oPRlDTqfPt/BMYTvmX7a6oZtgN
6mzc+6NTLFS2YVn456DBZ/kQCSOp+jG6AR6+e0WOTAfOn+OLk3ipwsJFFeVomG9102V6r8k/OFJO
BRrjDkRm8ipx4LI5xv7qDjJlSep+HmWhAo2y6aPz17vPPYxbQmZ90xmhmcSVplyvYUyWAve2Sc02
NIUoQVGZxCjiJmkeUi76+GiZLkN1SQ1dPTqyA4QTc8vmFmSuTjYJZoi5dBsGiMdh1P7xkb/K2D00
usN79uFBRoCa7ROMUnw/yxfA1HdxVjQh4tWgNki9DYRwQGp4oHiVcAEGUHaTzCf1bIllLZjAaInv
Yddb3Xj40/L+FTMf9zN4mVR90qftc38XkxNnEpB/7VSbeJKOVsRwS6bkcKb8BZVLRIWkdq+VhbxI
dat+YELxtW7LLpQQFihUdlUU01gQZqbIHjN+jsFAvsQCiJN0agXJCXn9gqBPth5kmjhFpAOzx2M5
LWaAdQ/01resvebnuNkWpkvDyiogJNFoKykgoWOlqKkxYIWqSealUwOYJgU6WDHRanFNDAglH9hJ
fTNiRZ8jv+ZCYP1eTb8Rl+/E6Ja9tIlKzR6R0iO6zPfyILnReSD3qYuRn3bVhktqWuizzXpAXKjS
jj3ybRoZD72xPZ6jx2J5bsX3ZNNA2zw0631JIw8TNH42S7VWKGf9QraRTGgr3iAN2WNYHSrfEphj
69kenQ6p4Uy1OLD8dHtvuVA9kBnSmRAnXZSYk7tpoUvMjxJ+L/vNH8ti1HCjT1fnC5CaMyRZPZtl
pOONyz97WFLTYQ6oVcORtHHMz5bDiY94ApSwuEyHSYqesvhJM5SAKRyLDngsEsV7PnUHrROdEw7h
muFvJnD/bebduqUiovgw2cJ9eyhr2uBxRY3nHaVpbA963i0VO6wPjaeteJWUh7fZYtAwmAjVxBGJ
NeHNcZmZVX4OTaILP0qWMv08mPt9m098Pd6gBY6ZOQxO7douAEMY+GKF9aK8ow/KDsZOFVOWf2sC
fPvLWSKHGEMhxDj63i3Bgwx5F8XOmt1Outs2+TGPh6eZeGV/AChC20NZhs1MLhRhhqw8641A1UgZ
7K0swASvvYiFlnfEVEKMzQ13ZtZUIPa0KxMnT+MI8TlgYFf7deEzL8A/BmD2pO/N3oVxpdrUwllc
BaVQh2fZftsiW5SVBWcxA63CbyJlLzW1ZaZByyG/V714vAXNFOtxGJlW8ofi3QRBwIZ9Law4DEKm
rCHiMawdtZWUxCJBOLneA6TjksQZwHxrcvLT1oacZoI03NkkOgfrEix4gX0cJr/Dkkuk6E6JAeMY
N1gBKdQpEoG2Efh+YxZlyGlZWb2Jv49sQfdSZpzqb4SavBgEKdyT7NEoEsp0zSnrerVol+dOqFeP
AmbbwRfY22kEC01CAjyjqNBoRqjQcnRT+iruwyN47TanYXBf9L6TcktmcE56lpxSIS2YHAuz51XB
USZ5dvhbO+ZcYfs3N4Ho+slsDRY6rwfS8p4Xf8uxV+PNDo7c5yKMmDNDID+1xsrSnoXxwRAXX3So
U/nFVQVVqWo8/R2rHkt/iW9mKRVe9DYUJAzj+VUSQdQplQ9gVmKKJFosT9neGu+/H9InrdvrT6eq
7b99Uk2t9Ng5B/0dZBxclzanSXO7bX1d2gBp5Tp3CbTHevZHTLIDB2NFY1LSxlq+tHGgM4sUisCe
O5meOKFHUphAXcwliORiVM2Bu5chhVXun0OMVKZ1n5OKnf0c34EPSVXNRw+bPZ2UNtxY6W0nM+d+
3tpzLZg7TmyoYWzclGyMH4Twdx1BtbzaijNObP5mQ2Tmz56gr8kGmQitDPoc3w1AR5d9Rk3y/AIG
FV29lmiI85Olnv5qcCWdmBsJUKmiTnzGw6C47CKEclsLXVcBj9PL4jDBiZfRbt/GAv2DROuDGriB
svXKkDiRhtpws1/6LLSsEyZ0Fs4oUyTBXN9mIefV02k2AZk5WbwYAbEPJwtYVpt/APIbGPnVRE/v
hHm7uRNv+P2w2NEE70I8KrhTBJKxqemybpzX/PbAtXTOYxuq4UtRNpKGsOeA/Ge1myctd4Wqm2mD
CB4UQTycdCVfUBjyNLKo9uzWDoHdEhsZTrBb5z3ejM9iNoeppLK33thKsxfiWhqYWPquamjw7ozO
1ND9DdaNd+DHvtWu09P3YhHaUUPMCUGzL7AgGB4syVg3f3ePQgZnZZHRRtFIjYEj0Rz1g+++mvnP
16FFNVkPV69ffzCH4pzycgWVbLaiFskcKWULHYJbR3uolADUIi0GYGNhW1omAB7IcNU1wiunVwro
Lg02NN0Nb/X0UnFtU4slq3PTJlK1gk3xRGyL1VrykSN/U5ipbs9Sxs+QmZFQH1ugySk8Ba0oHkqQ
F/CeDsRk5MX3MpsM7SmPcoCJ9yR18fGipZkdOhpgQT4BfwrshribHa1lZah+/paPZ7O8beg4PE5G
MQooKCITYxJ0L5/AsP9WIKf8xbtwPQGFaLGqsgo5BuDINAlLrsoSF9YQXlTPoKqb6y7onOZW+zvp
ByftQTqYjRv2yODLxaTcRDVMYOshMhxk8VggZmT0gByd4ZxmeTu+wtzdhLkqYeMsddK5F4/OdO+s
rXJAER+VlR91ziU+7gls8znw0cjEnpq73X6GeLP4/g3ZQcj060nCxwLnCvBOIZMtA1vK1bPbrr9D
0KYVaOsobN//VlkA6sdrNpYjW3gtkw6IbsjtprwHq9F7EyWey1ZbMJsYXnV+xbe0cEZtycZ3cHmT
OXzNu+b4p9x6e2xUDRV+H+QCIm4qmO/pvF9dg8Jnwx2Lrwi53mC6RiT6PhteUYVJiP0o+4LWt4Mi
/lD+YpSeMjO3HYiNoogddmzazMlLs9YAe3roNc66W5pZ6bR8B+e0z2+Mxzmaw50v99JTu8Q6FeF2
WvNutm0ww9zG6Whq3HagW2lRx+C0mu4rfK1XA/AHpmAfPIo1zKCs4zAXHkHXZKRLp5LOIuL094YH
Jhg3wA/g8/dpbreaBk5knNLq0mifu+aFUBnNmpppGXXNJdTC9pKkD+HKwdeY78vTnVLkmctf2v4y
uBObOYj8DeWX+uoWox3CsZ4vIYXih1NrviyQlTcR1Clh8w2Q6Vci639TSYhpM+rrbOSDlikRTaM+
3AXhdPuPOuRVrulBsT+3tTI/wDaabbF6el4fzKNiQbsPI0yvC6RqtugkjooKypTzpG7KPkH0Uaxz
YcN0GEyLCwDCBDXztTddh0GXDZMdX9rnYNpqLKtgdzyRIeYZaS7dqnVtBxcuQs+J3wBjQ4/6eXmk
Th257NpUOm/ZGlGLXxGS/pCVk5FreRmRkTj+KD1RMKjwx/ByRAeAdjgvLI5Oegj7QMrlkTRO9hyH
GuMa9RwHYrho829SYZ84wi7nEmN0rylzvMk49ZXYXh3hy23NlTTL3KkxTAXWfj957D6+L3vMcKn6
uM1wwhqZOzqwWlQn9uPPIMBYsKwYUP8fPEtd2eQYjB3Mia+O05icrrqXCiZ6tJ0j5CLyuR3ty/bU
RZMNgEnq1bh6pq+FCGwXw3To5JZf9PUppzxDgli0cWtiRJR8CFZVGBsXuJSE33jphJ9frphJMiom
hkznBezSsP4BzUbfXiQuslo10PhHbdh3/3mzfU7GyXn5cO0ILN590wPPgW20XVD6JRPMfwr5tdr4
TpP8XVH+53+f0b+TJiD6nQDHXVU4Q55oXeJHRC5QtW+Pw3tDh2Q9McVkrrcmbPpnHAg1aon913Qc
Xc0ZRpw6O3jHx50jSHJr+SIaiDHU5yJGWhM5k9pMjzxXcUa1iMF+L43HJm2PYXPPd5RKP+GATF7U
Y/FCZia5xrUJaFbbOOV19O2NZZ4VPNFftlKHieFfgN90mGWsOxu7MNebQZNLsyaPg6iglRTChjc/
KNo4qrsMNnv4ff+tWa8QMdJXGuj4EZjpx/NyUYf3uuLfntb1qYWFLlVSiWiK1yj+DrnLUonHOqhe
H83It3qceqUAtkMnaf9vcMveVHaPwR58753cNT9T5PO6Tl5YYQCuCxFAS7OQNnlEJOIaO2CSVNBW
eSV+XskLCma1x0gPdI2aHYAQfDiwziGStEKAe4dRtVBDlX5Z4PLLNJLOz4SxVTX+iXhfeYjv7jvd
oZElhMXKQtFLIZw/iheFnrMVMBXTHx22T60fJLobC+nIDGldnpL1oU8VbZi3vKQeV7YUGuRv7Oro
t+jgY8GR1AAduVGWlsygmHadlWsI2wOpfSh2zbTgr6o8PX/iStzOSXu0KCw044e6fo8XeM4A4Ki/
vKV/Qxh2DYUkyv1fQR8t3SknzBVIQBMauqxc76r7HqDV+r9Msg1AQeNf1ENw6Pst/Ds0+6nR0he8
jIGB+sURIwX+74lkcsWEqFo9wckHfK5PHQ5isgC3Vn1f6trxe6WoqNqwwhQ9XW8Azo6DZbSOW85L
Ne1NudLjrcA88IeyuLHeHG9CToMEWBxNrS7bDept4TDe4og2vNA0VDlfW2h2W7/+eUOaugOHjmpp
yPxbPYIINwR1VLbuY4h/LWpYdlDGbEwjjywZSfjHOSwaKZyhJTaFV54tIpJd4av2iL8lN9sYrA1u
vlRLROnV31TjU/EQ9X23wMQFx3ZB4R4/xVF3WR0HxJ26JpwWu1PDOddVTKN39GTgSjkHilJLo13h
0u6URe263kcH9PYEyRXCqf9TSSXPWkxkA4eSbeqCS4FScAV3/AfZi2jDEir4paxcVl/Qyt/1rTm+
Xwa+H1b1SJdHHDXr+KKEAno+Z1eOnbEXW58Wlz39g0tcwAyM/iStBhpE6O8FSOuowchZ7No4cAG9
1YU2QuPOwpsREcpnIj18lyu9qTCaT4T502YZ3CiyxP6o3dWVir/OaIk3FY8KFazhDkC1SmrRfsMk
K1MqNKy6+OkXOB8YfBq63+1UFoT+fnxp8HygZD2dRtLPLrzKDMBcyYCcxLtJocqFBsRj9+HEQRoC
cZfwckraopQYSqofi46TitCOYEUDE0SiG/SyfRE0RwNKpl+RtfY/N0ZapDKt5iXLXGsqmJlse3xz
ZNtVjMlbqMXEolmkecAmGqJvV+ig4OqI0vyITqtRmgYaBSyhTY2qdMvn4tjKh3mSUoJbGO7/822N
tItReYkWjvZ6h9/JPhc2i8TfgWothwXJ10uHUnPTpT8jpTmXvqT+m79Fh9M9yVw9szCupN+rbZkT
i8F+oU0HE7Vdm/fovLcVzUh3STV9ERMnZMGzalsJSj7gkYqamJVz+qHT1LhZCr2e7wwvujAEvhQr
cSdq+PWLZKfXmhz7CxtWxWjVRvewMseMd4p9QCYzVv4BoIoG4OO3XpBDjIqTCBuOf4WgBb9AbiEJ
o9WIAJGpcMnkkWsOgI92h2mx/Z7NNM4f9QlsOduowGZPizOo6dXWS/1svTnwN78VT0y7XaZ1fEiH
PFfPjD7Cz/nyajXH7/8mrWV9guLRqMuY2JnqdoWxA9Qx9X0WNsIlK1a8QW8kHQxMVrMSmUnwcWRT
w0SutwMUH4k5J4ahviN+rf41ugtxbh4cWeerbBLBs8EiByuhqfSULCOKdMUCh5Vh138J6zRY1+8N
zNUpzpC+VyRuq85+EugVTjS0+aCAcB82DtxJxLOzHZvdfAOSbO6qHzq0zV8LF6iddWj1/Jk7BhZh
MPKmttC71lJ0chg3FGR1cjt/ubzWcPn9NYa0qg5/q/Vip40Mjzr2hj6SBqyczMOrVBUWUChKN4xq
M9Wm0kwIVaTBlQ0t0SGtY1NevDXbwzY8BRV4JnWhBlfPP4txHmeKXijvjYd9XrhRiVPrbYMEDPxF
74xOTUiFwVF0RBP1WzDqRZpSxcEybOBr5Roz74DEKntaO1szEeszvohW9J77I81wWwm+G9df2PqF
PLFw1CqhR29DqyFBQyhgG2FY9jCvL+h9k81+u8pq2KtJbF+QOsENKOplcYe0qxNv5bS6JOFTtGd+
2AKD1BRnwksYoOv7swE88olGOgMoShK7n/3kHnwlcVhcPO2iJyeRTcEjE+ojwunpr8Sg2LLakXkr
nhjGpxjeZZhX/0eC+N09hvJNe8RGO/mZLCPz3bXFyQYJ9fpR1RxxeZ7b+z4GdBNqVnuHbFkfAV43
cXoGVKcGTMCII5BqDW6/CNXPrIdem+Tc0ooVnrq4F/UO/mVSLtWCfEDpfTBBIPuCqNwy3pUDlS7n
29MWqGZy/i3Xu80KA//nnCO+kyHyoLZWNzKG0Q1Awy/HJKwj6Q9F0JW534GMwBWw5BrYpnFLbeGX
YbZmfibKnKe/itNgVrUTic9WguOaz554LXPWuLElSnHkguofMxgM32SN48c7XT4DVYKf4BeETJSA
xGytqq+wEpz4dev2yv9wDMTlBgJskmJ0k8/xVd/DiYR3SgUExN2e6ndAx6e0clviaC8V01nMnhAw
G2dahN88gDzYeDjsjcxfM3S6LWUQN1rK3o7Ab0co/6pQn9+MNx2MXaRoMl/RwM5suYPlqfCdO5xu
EFP9ZV8viArjpW9w9UsuwhK/JkGv/YWgUiQgsOYazKf6oCWNq34e0ffgHAm4OCk9s7F4/5rC6qVz
+XjCtl5Yuofhp1lvpEEBU8tQ3u4NjitaUA72v2UAj5XQykhJickUl5mGySkjEwvnE1lCQ7lY2blQ
8KPhM2yl8TlNuquZz+Oy7Fg3P1Tx/AfGXAgqVk/zESoj01vHuhflyLsJHls/CWpaOWaTPBe4C87j
/cGtbmVablBkkDZ9H9A5eigxyC9G1z5inF9Ces409W2CAf2E8mEoLQ0ytvho9shMnRF70scJAQmk
46UmyVQp0vWsmI4kgq4Gi8URpJZ/0axDu/A+6bxvb//G+MOXTRlKcAyNMsdICeJGZqlt2Y0CDTzW
4EKgoeRVt9TYfeZ7CIcBGw3mZ9vJRZV2MRNIFLaSkYziFq91MCGOcJYwh2S3d7MRJDerllIrHO2v
H4DVJOseePb80ke5h94qadQOrjFjpGQaIkhrqBMvLnfiaS4bzGLPBxsyRHN5yrxb6tT4wPrXUVLu
Xp38n9Z8nFTsGYAqgFDySiO4oo7EHqxzN3iR+Q8s+Gj3buXQXJsZ6V7HvKpfBpRZb+0xrDxsgGkY
b9ZaMQyCCBSBCoz1PjsF9yF6fXDG4dRS8FSl27zoQIinr6DrDZHRwGXTA98CQwg62M2GRk2fCyPr
IjLCJwg/hs5qYSUvWflnBvnTCyqm5OSvm5nOHpaPEH0UEGNvhmALKq/cD9+ww+mxgZ1Oneo2iT87
t0NyF1CrKIEipiof20aYPXfm9/3MesvCBWe2+Qbe8emhR/GWcu6pIjZy9Zd7vJc5tDxHoW2q4lPK
zw6QNBeTMm3nx6d6TUtTSDbSRsPTaPe5zBQOrwTbPsu2Z/NmJojzO3CqI1qTaHN565kt3rn/fSvZ
eOPzGlvC5JvRTg/5le4nk1Lv4SizJzA//258lCjon8FAq+pDR8QXkQHWcTvnSTSMmHFyNHcSW9z4
/2DpsVnqgverqm0w1qFjRFkERG2kkPdrqLhznTHQamhdv18Q/YRFs98+T2hRDPggy2cQCESiBu9k
LkiWq7MtOx9Y89n2Ximf+Iw5Q2iN3PRli3mkCVd5KmV589BjWeiZhW3gdlqFCvaRVdXCEXqGYrby
2kUbEUaK93GYdDwOu9o85LPjRACjapQYLUSGXOCZVmF1ewMQLWqSuQS6eF8SOm4ZCYKKcHFfOj/e
ddpNPosWD83LZCzQgSOBpPNe4fYfvjK9iebJ2oj/JioJClNaym/Yz/aqw6D8SniKrd8yC9MWQyhG
AyFwT0HXqyZO42W1f9X3EPtafXQayfUorRMiWXfY9Geyo7YAGDrlQ5g2y++4Z7qZnT9PSsOcI5/G
ZdPdJ3ikiHJ5lfq6qHJP4HT15hPU1xwCgYU7+VquXli1KOQK6GzY/WnbSb0q/YfGqrJeTCm7SqJ3
DRo6dTOhRMqRz9y8fL8GRFCTGPVj1glxKe1Cj7+83TO8HgfEJE6sGUI2vhi/As1SiGcKWsV/T5hB
VtF6cc02QHZs7W4+DfynWSf73hkJZ8jEKaHMtn6mG49HoCmoxdYim1OoCpqL985UjP+82NUvorla
UNVwM6uvRoFBPBdjCMoe4ubtZfFfvoTJ3W1HEKvbztYvZmbnxLSex8nXMJ5gol/OnS2vrV55Ksrg
x2YoXGuYbkGRb7Ej4yd3mMAEdJRIWQfmS95o5NGNTbEXkcju+p/Pi/9re7S60JcUzhDjXUiYWBuB
c0PKYg+MNR139HA+6fFMgQT7EEqHTO2EsiYKiqTB71CnBLR+fKoyM2TqI5T0GT90U83eF/Rz1+DP
bYSsvQhCkIkloaCLuSc5j7aak3NMtoEhSGTYspVRajPthSPK9SqTbX24ntq4Sn8mcfp7rfCpIiWK
fe4cVpR5wAn2s+wO+JHwFXbmn6c7ncgxtj2LgKzrXKnYuDToQiX0d+TArDlfk7Qg8Ro7wFwmoeOf
VLnStAhVANQe/5AaqazusRfw4BDgiPrhaaeQL97wnYtIG0yIcl522vn75zQugdcNXn7LrKlZzRyH
uhEq/KzxAWsCt6IXK0Cta/CPV35wir0Ql0JRp1pJx/mfhCLZU1X5rmmv7KTX6eOr0qrN1sUfL0QU
Ge9iMGRe8xByp6v77Zlrj7KiSEEyflQbzlr6aJnlEeonS2JA711XcNdY27AMs7qmsKqIpFAVlI5F
kMF9qvko4XZ6zSYSWJBh9HeEuU8v+dewDb/pPxiJzJBRSURnuyc7OKigR9Q04Bv77WF4yYBbRjzS
TzNaa/es8OsMG4mMBUvAjVg7qwp3huHmQF57xrnVhLnylEeE8QO4j2mJxd2ZLpWIldJBgWvfqKx/
B258dtmz6hLFE8i+5Rukq9qtBlcXQOVpCkQFMlQk994xuKzrr/t/xOzhEmFbA1a7ReT/d3ppIRLJ
bXijektxoqBkb86uo3mao1PK+KZ679BqRbzya2q/HcdsPW48MNr0iee4t4Htru0Fuo8GC17NQdbw
KaZK2G8orU4mdrhGQUpn7eUHPmzvFMB39WRXvRGeutSWSCLPfAuZuPjTAbrWEbWrD7OjXdyrVhg3
YfYKwUn9JIIfvRX2nA3YMzdQCEG/MHnkejESoK8GkAEv0QDAQebxB1yYKig/cm3gF2lNgvlUqF6n
1t2PLN84vz70OHZxFm3fwaFXJIEgp/CAlK6Ja0CmEEGWgEJGL7CQqhujaYXmBJWjnB1LDbgkhQU+
RnbGt8wS3t8Z24BD9BqiLoCWgVgWLf1HNcg3Uxahd6So2xmmvX2L3k064OLlVJgkRX+noUZcwdon
lv1+f1IBbtdMoZQ0hOs413N9fvcR/sLBpgvsLAmgZCRBJ+oW6tPuDQRFu1Z+/ak2g+WRsuialEky
WXPuKPZxq9Ju7SSoNrdUWYcomaucK2TaQHnzG8HT2xpkesxIVrbRR79qfhSX1e2LMJyaV+duwDd/
Vdctx4Vf/1gRzyE25S7in8s12T7RRnQ/tUL6r+MT/6rRaCD9yyEwFqCuRByQ/V3FYdywzeMTpMY6
dVIopQUQD0DfCIYBf2ml3iYfcF7Oq55jhYw+p54xo697F6C0ou99nYKgwBF5Z8QTOU8iCuwyXVQC
sWiehoEMHWKNMKUQoX0hnQop0Q52jftKSeGrTP++hmIxp+OpWUI7HyVwForWpLLdyrJi//kwlnD6
h51mS2MGbxguIszw9Wk5UTfn9SDfRGWtP4XyFArDTsZ817ExNEIYQdVJRk2ZseJ3RqIV79tiokr8
dtE/HBJxo6moQ5X1hCgOWmfBPimMAMGlqPFdltazQ3BHNqFXePtmQKi/dWDKbkzPTe/NDbiT1jXQ
htPkZyofzmTbMs8BuHIVa3FUM/jRg9v4yUzCMzPJMClZi+YqmKXBPLrJnIQU5Vy8ajz8Y0/iMCYA
yy/CZ1MlCvw04fz7ENS5FIEWFsHBQ7rhqIdcSVcCR1fhDP/HKummvAe/a+5eLBnJNP8p3zQJNg6J
L40OsubQyFom1TxovueSy3r1cGrz+npILpPL5fe9ZCQ89Z9kuGao4eP7GbkCbs0idXFU8YWvq+ST
Ch1gVsIXUQ9yc+T/598+RtrG7wtA41z8b+kShwfjIiKcgarujiM3qS9bvT6UaJBAc+l2S+7xHLF+
UfuP5MaKfdQln8X1xP48rVoihgFhLTdolzJQyHVpuBP2Q6Uzx8+OEjB/zZLeeN3sbUkWTIhAx6vx
ucvx0Y80qnNXPt3ZVgApt4ykKZdM0o97ivZf0dXQNFD+XJXgqvclRlvJLHQ5ZmgVahpIEMCReRMP
4yfL1/H+zRoP0MZ3AzW1WOUYr1smG4JtXL5+FC6+NfwOB2FvhNMGsASqN0/K8FGUtGy4q1mD3MbR
RLWh0jldVOkWvON04ugh2fvlhmYTwh+Yael4o0k/no6hfy+rbQaKPuJcU8LlQivW7uEWg0Whk7UB
dmWKsJhNtprQCh/qTOB6/Vw3E9MkOlwT23XU8vjbUwDCrT+dAK5o0Oz6gXAP5vdU4mPnzWLdzanw
LjQD01JyHcNfBuSgPuMpPYQ+IyFZ3/Dt34f0kNk9xV9TdY0+En5UECJ9vPXgZMl3JnVQ8sogjeZM
2XZ1bh5Ij0N7dpvOgGj24Tg7v0wS/vlQMYf77kv7CYm4gcSQ5PfI1p8oLGksCDFHU6iYFLYpLOQX
81j+XhXbmq4c4x6fBagRLjOsgxadAp1o5LUcSY1u/HWL3ncoz0aylk/a09/O1d//k/++k/aSDLkS
o8tt5QN+ROGermWOiYP2BA6wpZDksnCPal/ukr7GN07mOXeoep8Nr2q+jDaliBFLg2nwIuq/sKMt
MyiqnwCVROFPK2YuwVBrpDhz1Oz1AqmuQED35RRn0zxzYPjl657pF1c09jgJqvv3FNlnTMjtBtpR
f2CBolBQ85A1rlydu2/4XNrCx5w/+OpAy7Iuio1YHvHzcaq/dopL740zBEeTdxLAa+FeAOF0SOrS
i8VpJbVr2ZEbALm5oIicCJaHsQ1MZ/AQzgMORAAKFoJr0FFqyIg/hdNnh8COI42WxVcgxKysc4ou
/yyxvuj93bWIQ1q34urywhh3gpMNUiONgxOVrO5Wqahsy99E1pMQKG20OQUkZHw2wB6XnAFx/gcz
CbEfuM1KDSYNca5/jEsRzSM+yjeXpBJcaqu3fgPI0YweImHkQuIuNch+vkNYCMSunnKMj3gnBYPz
qNJ1EL4ncbFRdF87EsG/p1aPW/Q11Nbeimqt9Js1uZk+r9k+IPcfc+dd0+e8WtztNIgPwZTer0ku
TaNpsqucyydpiJtaaHS9lEkfzX85s2851qpResvzdemIGWSjjgo4F+qczEhauNJ6lgdz1L7YXbRz
t8GCOYPVQwGwDbI7KZaswk6RKnLmXsKP+TZqIHjkCafo+bjvNZrxq0n2og0+C6XDOIWIPKziWe/h
GH8VmboOnab5V70X1D/9n79I45Oiss/2YhmDGk6DFrWibjnqqQgXOPuchgTu/QTMlRLKqeAPi76p
bt9fRzzKGtv1G3skKf4HXEFU+CNaB1uZNQjPSt4cr9AZ275fwd9PS30TVxAWu+d09HeaPCZK3vgQ
iFpCMoT/ZctchowusjgwjpJm5qEoSy7IUEI+I/8SnkEzLecwm4/N4a5CZa0dOkS61EnkFV/sRpkV
BrFzt5YjdHaMtdyVSEkZwYtDPwPdouXsdzPTn9iYR0kiY477GuqJubI3Hw7mCDYNpCqhJzzxv0KW
bPXiSDiKykvgEEFLdEkcubFflS9IyGdKM29zTzYunpWKfS8HfJptKa0zPp4nVroEJvjradTi89WS
/mn3io9+zanZfVej1A4EhHb1UK9SVcWp6X7foKOXuI3latk+TwZgy7zkiP9pSLoR/io6GmAV3J85
8qw33m8P/p8yNWK+wfJm0o5jxefBls8zOA7wBc+enNVUqe8JrYD0DAUtecpaEynNyCBFHwLpPqK6
HvVPGTL+EDM2SCRp+8T+PtKXw1zYcGlIqLvRVSxp6vuVlIpNpkt2/MdouTW1ic+3klV7m2US6Mad
yC1E3unzA58QUEESw6h65/mncVwlmXh38FhV7p4WyBk1h6SdLIghLIl2A2wXO5W7eFpVFYIm1yyw
ZCtpB+DAPjEwhxyEzgmxX9dHYktVo/K78Q4cPZbZwATpYTOpnS14vknApCb8pXd2xB5zN2WLFv+U
caNR0ixa8Or2UPzOaD/gGMNPvdaNdqo3hTx1B/BFn7ZEhoKeRMGC6gkWwtQe+AElE9hYtXo6qkDi
1t3OG5kkNCYJxFQVmMsr+YLeBxo5sSltTes/+ui6nyiFdUurDXfIFovOnwa6OYe7Ytbl4iDeJA4d
KUYipXcoj+OYFI6Z5R85OElymVNtNbc2gxuuzdPfQH79TDxSEMwsNPRjOoP9W2F1QUe28Su8TKP6
7yX6GGt99G045qCWlpVKMRaqIuEqeWWmCsHCC3tafud8An0/HYwBGv5Q15EsKeqg7IqlMKQdFy/u
G9XeJb++GTVdg7p+GmqM6qUZklFNbJMmSfahgVAInK1VI+edKtp3LetvAWc3WlBsxPruSPNtkDbR
Qszyv+i7Ag4vOCjxQU2vKI81pMDe9ntk1fPUt6BMIG0jfwU5R1JdwzW59f7u4c4PWuxFUojXOzns
mphBxqsh5ZB7OJ0gQQRM9ZdNlsjfTI8q1j2Sx6hAicM13kB7Fk1zlj8IvZP1VXWXTtscHuhDlXk7
ub4yWV8KYwwEo4M30jfhRznrO9uoPUgMHUUXkQsh2k9yiOTWPTe/1EotLCQpeEcMqHPerIP63ERN
yWYol3PT+DJ5QF7spIQ0qDLeuioQ2b8Ha/TeXtZZep2YkNtqFXror+k7CkCNpUpJ2sxtpkhvzJ4S
H8CKv9Y93twowkQj69PyuZu9rMrMCmNzDx5JLMczEIZwIGkoScYfv99hD7tayrewVnOfHQfPqFBV
p2xRw3KdZ85jBfKBgCLGQuCv3DjdsEftzOd+Y0rW8gBKtzNC6jWuLGhcu0krHbMa4M7DwWMWE6C/
w2Hp1x9LO0xqIKqcE8l6Ipqonp8GgR3tHDzG4DWIo2uBXP8td2kUqvpPcgw1QnVFWrRe6hDNjUNe
StO6uwNTVX0lF0d3r12becKJxt9HwsxoBnG5v+woNobtUdxYEnkFGZO0voWjydTmJZd82xUDCDop
Iviy/3yosPEfL5z7JSt688B1VIGZ3GuwVm/srTONqH5Ir1DmHJmX0HIHOPrWFhi+a3y8LW7PQ/Fn
J0TI/LzyLqTGrlpZida/yAn/nGoDhpf4w/+KbrsqOtYHaWfROz+M6Xr7WJhCytsIvlpG5qyYxchr
s2AC/afDCjPzxips+H+BX6sqagX5iycnwTJzmbBBA0gH/16ly3nPMzeGOcwLDtq59nWQ8muTQ+gs
0WpgHJsxItJ9XuJc8BUZ6NqBeIG/MAzddoDL11ve9B4AZXliKULNM74eXvcwGm9Yx4GOnk6CPjpU
OXDfb8c09XRCkVpjfhOEHOfthRaUa6UE6FBwxH8LGZlD8GdB2ViAO+k0CNgKUdNV/sppD+GoJsl/
l0E8+qL+pcgo5DCdtwDmNkYrJWjgYNHaL78FI5/vZBWRuLdhQJE9RXcMwMIJLdGGko9hAc/LCGSA
icW6TSR92oOiM4gcLcsIAMK2UuGDaYwImFCQE/b1liDaWk4XqQYdQ7flAtzDYGTV08+O2dyIuIqP
iVBV2z/Y63xIm5RtnWrs/tH9YFBaqZQwYe88tdR6c9GvvpH2XYOB5zdciQ3TMXGRpcLVJNkFq77j
DwT/K++OlGC7re5zu82Km9+E6BT3zmHT0+YKIWyRsxowqaYzd+YVd9mQRLW9qwF05I6X63YrAZkR
ZmeqlkdkD2dEZH1kSc6aPHkWfxlSvL4rWAx6BHjLAv89FyORO41Dke01jRiUcsTeodtZDpJTs+mM
gYL21gzQMPrP4CM/iSsi7KftC5KfKE+8wN93iS6HGN5KxDeGbypaJ7cIRUbfngCzcbmQCn9vUmhp
8/sqYCSg+o2rgP0Lc89uCeewoKYKocx8Slh71R82A1PliVmYkswLZdGJ5dI16iU+ooSrKyFjryLx
FAApNdDhP6m0JLl1V4TWAdOJCLWntZtZcX7SYB18/DhNnEdWX+L50r0RjkrRKMNX1C4h/qNf7c2f
AmfpFvCwr0kQUdB8jojqaFoJb7MBcRPjjvnkmOJjpz8ItkWuAQ1xpjfvNFugfY09OWRYpXYY7Fe1
h0I9LdtYUQ5Uuo9HiBLlFl/vlL1zuFaVYpHSAuT4mswmOD0lzinnvafUGu3xOUQ0Vpn/1i0BQ1Lm
Kg97p17beB5jHOZPY8kKo0VBeoiyOCrZVb78LzjtrET2qFOjZeP35gGBun+gbOH7UPD3/FkHXt8Q
R5WUEptZ76ioahNbf9pDRpIi+eGROsb91/eDqGBzBkXoJq0/gXxaXiDuCtdRtAvzIiDl8hsCHxvT
ZFYAmkhTq+5nxA9a5RCPfW7GbNZRQgTaVZoG+0l5j3rAzX8nI9SrjYQsdVFJhckNpr3v7IXG7xi6
Takkc7NHbiEQWxrOXO6dsE4NOS/GBwxLGlbyMP+u9OnosEzFRy43CKk0tVfv3kBRpqnVAFl4iHU0
t68AcgBuCant8FnG3Unkh5lT9J8rUmfHKzIk88gld1ZbBoEM2j5EZRcQGoz8wqra3Qagpz0KogkX
E+tKQlG64sw9bIExi1T6T7g21ZI99vnDpu+6BiaHxJNHe+dQB3k8wqIf00upeuqFwmYJ4KF0eb9N
qaspAYAXT9Jg1lFklnvIQsWd+tyvW0aAog5+VqEYx6DepXCI9Vlyh1uM3/cbAq4qJ1Jg7lYJ4cqm
OQoMQmmSbvzLt7G/D97L7x0i7L50Fk9uMg+99r5Fk1WRzO088v9bjhTaCeZsDcqHeOGnxc1VGjEX
TWSHXWLS+E3E/FV6W7xIAwqW8lf8DGP+XUwUG/m19BvX39gNS7hIM6K16RTPFicMX0oksFe+b8zL
OpfphTmT2Ry2MWSzW7k2b6DGMwdeX/COMG7E5vjdQ4EyT5hu/quoXWt7z7k6LZAsPzk38BamG3N4
llytcvIdwbwscdOWDgJfUdfrkhqskuXaSQiAqdv99NSei7zlRtPbYiboB1eL3WA26wkg9oKJaSdj
2muTEAl6jiS7YhkXl8RrwvuYypz6HbACAKUqlV68kIexlp7/FpWfXCaz4+YxAqskO00oSuDKLFnc
ryJIfQ+Qtq7omUGs8Gbo+JQ2ZMYWhFk6Ip0i3CG/fQv6tv9V58PfEzS/KC68C1OgHh4lTV1cDfSl
cPHQ0ZTl+Cwvbq61PQxrwXRjeLAsJaDWH/0e2GKKFZK9IeyUBDWzIxM9soZlOb0bWWpjPsJKt5U1
KNi/1x7uM6wIBv4ESyxafwJN+0GRDCk12A6ptp8nXnLjmsko4LiQVD5vLPpImmt1C505zV9F+jr/
CxPg3mnlJYp2xLzAfL+qaTXNwWrxRSuBMkHe70bWeMe1CQWjeUR/m17cJxcTRlIPI4zxPrd98dXZ
T4O4fLmRTHACeHpRdUSFDLEdo2Q0D3xVXoaZGebDRqD+ZlgBh/2bB8PactF4HP++2q3v8BcLE1fo
fuIRA11kciYUFEEFUvl7J+lh6GE8noWzHh34eYJjjdmiNfUsayt50b5DQfm553PcNCvJ3Z2M0urE
vYtiKqazHFAzIbbwhKTVPGMTrjaVqxOw5iGtiE4NXhAL4jBqAUa0/VhCQVmKd2SP7NZq06Lq1kID
F53StM48nalp3tai8GGLzs54lC0wyGdMu5d6Re1NOVdEXUVyT/ngwJDpGZO8X5CbuQzYu2wSt7Gv
S6YINKV8D8JQkghURjXW2S1UjwH3wyGehQe+xk4RpYwztGiIHCMPlibDeBDaHWkVFULTu3fHcOIE
9oUvDO31sVKjc9SyAbOyMh6RN0RBxhhYJthfBqRgqXfg+pXVrd/Jo5DpubSVnhajaDaDdrdogX7r
71b52fCJCumdgLaJchzlZ8i99ccu/TuiHqvj8s7ymuo1c5/KqUm6JM/uSWWXhhR5nWZqXrVPuMA8
BpRsuvwv9aZ87chyrsgMyk1XnH5pvr6DQk9Xuuk4yQAy2AxITsVpxlTCPAxE0+nT0rHJeRNbicL0
f4wpPuOvX4GraHsLoTQAoah2kH89AVN8ncKpmHH8da4QIx8tGfCNB3ePbTt/Nx8UBzFJOao0bCZb
7MDMpNiksaC2FiPoJut51sPBcpFP48zsWapEC+yZQpQ4Bnjn4ax+WOmaU8Fkf7bAfGrRkwrzoS8N
VBnzhe9J0IBJssb8yFPcO3ZDjpJimNauyAzHlmPrOs4adiAtQJryghIJUPDlkayHFS5E++hVr0X+
dHR5lOo0rEtUVBc/aSkfVZRtAmvnJwpMc2mkPPSTkMGYylLINlXEs+LBlRch+tDRbk7jgx1m2HJr
enY3CCPrd6yx9NSvYAjt5psn1j2q0jmaQ09s5a1Yowl7464mzmQEdoBmE72k3hT6n/mZQVXUMrJ7
sTtsES2fpmnxu+i4mcw9owRJUaFNJj5zIFa8IY3kd2K9E5o7+eynMEeh+SxitvlC/IcPDdXn657t
wbMqbfk0wUbQyYLe9oLV2K5LUvc1NXA2R2bMNALUDe7B/p0n3olZGPJGxGpGgsVH/YFGdtiy63ol
nBVuJgTLOb9ptpsBUKlBonbsu44DFKpMCWtnFdEE2ZNOwt5MRJLrDvUtHfcsWHby4FXy4cP9pE55
jSjlGAAU10OELLTnUpWcCXrRPGTz/1QZ56OEJe2ZNl5AzeeAGA8TUvR3fb3SwaQLUlloVTdzAb0n
rCN/UwxXeTY+Cxhzu+0t05O5+07aipfdqXnNBrxFipd65MuUY3rQjFwxtq7DZSDQ+jzWeCldvUwM
yASb5q3I/JiHBbVPdWSHaVvrnEuq5NnOg40rlSjWUlADFe1mer965goVPLKVoOod6XDyJPhLdkjH
K7znT84E81cP6eN/YuuUz7N+AJ+iPRL/NB5vSuSabBiLh2Uv4KH+SfkVZ66Xd3oP/skcQVTzxN10
V2VuXQ3BhMTpVhYniCoBYnD26mUWeQP4XgS5qRgZYEshTHHpY3nUmYmAhafD81rKpKUxR/VW5T4y
feLxYUPLUFh8754pGmh7q66lrq18to6/SCrPKwwYvg2sSICeeGPTc5WnO5EXAqjNiq+d0wg90ueD
9Ik5Eu+ydTdpeGxIDXcxj4mWRJ6cYVxzhK8PR+IoINdyI5dtTUHIKO2430Ur2NZtkahu5bt/G/WY
7eQ2/BgIdnHknerG2NXbma0m3zUwWT8Nl2Terx5J0DRm9n507ig4Q7d8eBv3uP5dU6ukrQXkWvUG
tVqju5mCYsnoUAAsvgP/l3mdRhxdwHAq7hKwoQBorFWYqAdZvsW9RbMwMq5Z98HQofXlsZSpsizd
AlhW/tyMp4laTy0PvXjQsuGzt3SyjBTrMPZNSq93wvuZc0i2iE4kTWkRAWu+vf8zVY5+tdU8GMQT
tVRSc67rAKY9NesqLuG9nUiao/8eZDbXlqnmHK1Z0R25A0DMovkrDXAaLj8rXPcae0eoemoaFZoA
J3GEES9oZL23kM4YXp24Co0fEFb4AcBfZh9EAzTEgnjPMW7ae98D0YPE++F9ta0wInbgKyj1sKis
4DM9uGcQmrfWpAzfGZ8v+l/MINAyd/7Jol8NcdXBPI1gHDAzZfIOjVt1n56T3f8m4P/KO7QPwUd8
T8iNEtVKB7iq83BYkoWyF9BipYUQOdW0gpJYM41/qxuiD0LllQdrh85OR0JT/oG5e1u7OFZND5MN
xwioPMvORd+AkpJGg5T6oK60OXS93raIZXEZT97tIpPnuLxJ8FS2X9/IkLyqbOyTLflbBanoc+RP
2qtTJF+yxE1ypTwVlG9ewRXhLPohURGA92pzxszT6boTibBgwgm6UZG+EaYZ+IWNogpZ9hkudnB9
aRYXE/2L6mSjJp3rd76Z1s2hQoQMF3HMZC0b+dLquYMVGVI42n4yfxSdYQ06jFO8Hf31nmhv5I6p
orixBq2dkQXJIBBbMGLnfcrSw4MlZOghQ3QJ8D0gF5ZPIqfHMIVxEQXd/6KV5Wtay1vI5CiYnVUr
ebVkwdAmvFYgyi3YwmQvJEzs/ebw3Tr0FjZOxxrSKi5n6pxll9TtWrrFRmV7RZ6xTVbx/LYLLglY
tGGuFCDbpuKtzcYXSgl3mzwDTqIrtnYA5RR2+Z9R3Wjgbt3AV3/lsqFw1xpKTcngrm/2+3dVSyaW
OD9wKz5a/j8oKW7Md12nhDa/eRUfKpf6Dso0/23Q/YnAT9H0LlQ0q9tgYMSycqwIlCeo3ymlxfLw
IdxFh9i+x2/An0MFo9qTgrluDjIGfUtCnTkc4t9/QL+SK22U6b2lHhlNzPIqCUw3hah1TGhoYpNs
ru3r5/eSgSRuLoK3lOrN8mQ99PqXUVJ3IP66hu6tEcsdo+wDNejsEboViSxvYmmW5Hn/TwY7Fp3J
PwzbLmHsSFlAvctyRkskoyoIBXqkIyOGFA5HlCtKsu9/8HK/wxVFaoW5z7J6rY1Du53h/2eygKg8
mrcAzKX2vImdT35MB4+jx+iz5nnUVS8PFUZvRm7b0CXoKeQsIETyw0FQHu9JyriShjfMW8VrIAzR
RFd3S6iFvmVAkL7hY9aVl6g6wKkcL6Jft6fpDtxbKzgNLUXsH4dDJzxE1oYrUHt3PMqGX4uQWtNE
7m5usGOv/6zobUo+sxXnR0kAwwOCr6SK9XG8tc7DiXMxglcosRwci5zbLkZoABV2QsP0KfAwjNBI
86p9XLkrnPGY9j42Z0MUZulq830dcwtq4wNmCpX0EMeeOfO8iS7qFprhWqFm9Yc1mb6wbG1t5gYU
zuPvWv/g83CRmySfIICkIhGFEzleoFkb8T9CUD1AbWXM7GHqvL1abbptHQcOiqOEGIAy4BA8/Bzp
u/IHz+7RAOwOZjcwFSsUQil/amoxkubYn+pdMX4u4UxIJoG906XHahWAFiuDYU3Z5x+f4EGaEj/y
p/J0E0MRYoaNdFReKxHgbB9a0zR4sUW4DuTwcRfqrIWoeNmdRM7V+uX5FF2ndk4trIqQSBvxxW2q
oO3MBGQikH96bxfaySQSh7psvfl+kioTiX+D0TteCCVaEFx2Oxp7Mxeu0JaaaaokFBTNYTNJjfWB
rfLVKvNqz3fK1LkCT+vX1k9OGMkadfYVpSPUTtT5HOZ7trQAPyi0s3SvBgLjxAj62bRfBltFY4Ys
Q4epWn0H1MSXpvIUCuHs4QU9ONluHi2jxZRcuq1om4aP/n+aIymB1U7mmWP/aitqmc5aLMqFjQb2
bASjCEkXvk2+eU30u9KJFcEgqQEBN3mfNxlyfHr00yaHetWmxC6sQEizvyJeB92h4r/ZakcLtT3B
56uOz6QxeybcVH1ZzkHUIajknjlPaHvphJaOg+/5/D7jx15s4OfVhvgEG7iAxQy9ANdqAE+1ipx8
RFsCSV6i/HiUd6JSyV342UHFg36XrTHewovzEO1x8JTwQGQwznoY8kRl0kchOLi+SF9poVtX2+ac
LzTn7kjsq25KvDgQr6pN/DLRf+7mEjWPJBj35AbJrRIBu5LfvgwW1uR+pivPbENh0akJdSoUSV9a
yAyJI2ggxLASx6Pzc8n+oVqOZtn7Etg7cRJBNQkamUSP//bzLcb1WKGumfwF1v81jbjdlVBjRZfn
pjjiFF3Vwt/TgEYneZvHAo5hYhIsfIJ0gMu/A65yNggjH/qbzQphTKxgAIscMA56Epv1/ynY8j2O
YvlHmFs4UW6B2Y/TMHuGN1ACIJEhMFelU3ea4jeL5j74M7PY2FfeGLYdpO8OkojOxj+mqcYDLnEr
e/lvuIpqc/NohiAijX4wWFnG9rwNFw/2I9DnqIRyQgiaqBQTK/x3DuMI0t+X6kkR3Ev74W2qdz/9
0wmGTU/MOLXyZEpp5FpJfp8sFQAjpAhtE8vZkM/BSzRLLczcmGmVcrUgWdJlRznuRCav44EvODB+
hTnL+y4QddFOj3fR1ncJmmeUZERg/oMBWYyn777UXdeawfNIsPe1jooL2ObkWW0Rev5n/DHDkGs0
E2+NDMqzRB7DHN5EbPVMLkTkVwDJ4ZOSn6EkbY8BKUENOG+Qzt8/jK6k4oqBOfrOGXyZAWzR8j18
2OaNevD7U88lhoaDwhJpyPXqFymimGGgjLJA/JQkIe+uoPwKucHEVcb2y5X55eFqUDsWArtSCmyB
Yz9CJ8rczyRgi0F/8seyS7NEey+GySFXA1ytV+p6Cvo9CPafi2DAk6D7/PUtFb+ce1jhO3sikkFs
U8xKRdROF07z4ogJecbOitU//ezpwQSJcDiFoN4/BqoYHFRrN29d6Puaa/vhrBu8w4UcI4CptAx/
IRJRfazl9+yNuDzFAtQ0ESxe+3uWWQ6SSdocndP1AcgNBZ8IBgef6Rd1G3TL+mwoHFZ+nZGG18vV
0o38+ytEZIE1SMFWRpgzMnhDOmQOzUEXYKel3606+tgou10ODTXOHBQCxG3dickGHzl5NAXz1ROF
C1pOss2Ox/w/VPupZvJ4McGVPEcg4QC83rh0A4GZtSu+/QCJg9mzd2wT6PzFPP82Dv1xc8xV8vW3
/gkgXXmSk6f0BJXdF/kBHpWSE0bE2lZ3r+wVdY0vD7F9QNeKfZTE6BtmKwrsbN970o3N1BHdJ3DF
pPAo4Ek1jOVrzHl72qmBpsCvo/ZS6AF+VKVSmGn235gG0Sm4PVKpMwmsHE57EPEE8URcwXdrDl7U
FJCouY9KeDM5ivvfCPsajxuDMb1qugUJsLoTf0pZ8CgBT/uuZZswyyrig9uSXJihx/sSiFRsrpTV
CldaSEWC5aTV5ATScqX9Tsbu+hCL5UZbcj46MGakOnsbT/kzN5/G/RfAJloncHGnr5Y5TDYlqcge
mQDUWxzDg5MEzjOtgTm3XSmxWmFZXlaJivqwS3SnZJl8E4Cj8ZUzHqcYLPvy2b7f5lSVz9I4vMPb
7hOhHYkfjU1tw2j0SZtLBCCUQto4vtfq7PL3872lErylTuLQzqqM0zrwVAMumPjCafEQZqEDN+4f
Az8q0EeiacEBNd/DkZjFdhyQ9e5QSchMm3GQpj6HRX1RNwxceyRIO9wJCCaeDimz9F/sdCFZdGFq
MUMtZyixLqnIOquGX1GLjVDmEkzzkKf1vcXnNtHFB27NojwXmL4pAuFSi4ehTyGmmrD3f6qZlSnH
Fitkg3wyGHe1ICvVKyBID3mZh+3dwz0QKzp5AoTS4dsc8hdlSBQ77bJjC23knk/mKOzQGOFaJXMV
UjDN7F8LR6L+pJWNbWWTrwmn5Ecq8zOe2OJvR0vTz8S9APvnNbRhSj4HNETVXI+Iy63KiBiVvZ3j
Z4k/oN6+oZTIBj0ACdxa62YoLaFasjgAB8xCR5HhknkiZRnpTTc9o8V41DZ2e0zjkcAtmZIAJLEj
PylZV3YnT8wnKQPIu8qg1U+45UIlicf9NNPgA/wxhp6o/CsaoYeleYBevE04sJNaYlxih6wxAowM
6uGwpoDplWE3qQDwhnC/yhrSJ2eEUnpLfGIINi/cXIyUwarbxR2IecvTjjd0h4uut1velm0dNelP
U1xw2kLF8OViJDOM788wsFRk7pWXL+V6SEjzVUMQoKa5VFSCXYoLirCPmdKupmAc8J73yyu213EE
kTmpOxLeTFeqTran4GodVewFPVBsQegx7oFFN4CJyFhCBvOHpuyCRESjOcfduA9GmZSsWW5NxIdl
LFW1CMF8WE6sUTcTEoLqPE0ZXForEZ06z0ONlFHScfTd0iUHdncjabgtRFWUdTsMrFAQEeKc5zGG
+VC/AaxG126wck4CeZDuUGBNeR3UElWTdaM20+D8COQFrxaJIxGvP6z7T+99TDYVD3VsI+VfmgPd
E9voAMPnnb9hv0VrwUVlgAed8vmlRUQ05ul4xvUE9P/wsWIHhpOPqgcQ3QUFJAqH4HIKEl/Gfj9u
Wv+2nYM4TLiHNqqQ/hkWwigBN1W9vNPnApo4S26dybT8STjbe/SzJA/T1FrNgZyVLZ96j7NUpkJq
YQBToSiuen9acOXjjkRdPrCmpI7eP8AxI8Evw/Pe1bBGvbjY7c64F9ivP7haChD5YKepYbf2Tsth
tqL4ST4I5qFC+28UZ88knGarvYkvt6Tvt47jLXd6tJ15YEiOPNZW4yl/WHcpk0dtM1S+9iKTLiZu
B/yNe07h6Ozj+uUaLJzif57yNJtqzDFP1/sPpkqX8vSko+5QNGCbjZublHSEkoV+32whCL8/bBnY
Vfknkqx3lYylExANocW6ezSW0H30b0a8NIkbeMvnaCb8lqjoCF4uvDFAibf8cLV4ieZTyjEZ4QFE
srfXn6x0szqPY2N7x6Du0hgKaizObQ6sfUOVb8fDuzCEjRtEmKuJY3mNqXzz4pqt3LmmuiPaHCU9
oIAs7Rpdlo/BqkTyoZdwXIs8okpqplmeoB3RHtbpBm7WUIch6wgzNBtuQd4oqCvk6c+3GDAcGRI8
c9De8T1nQu0HvXXo5dsctyPVeiNfoBKZRglQYy6TziOd16w8zivgI1SMq2Z2gfAI2/fM2J+6dvbq
8aCBQf/JHZkZ4xDlK9lhoTBdZCZB8w2yr5CPxcKlQOuNnK2p9Hhf+0Lqnmg0eXWJConLlNPKoFxD
n1CYcJyL4PviQJQVplAxaWl7aZy5BtZwXy6DjP9qia92/U4uoWuDK/Q3+09PAh0ptgIA33zMBfa1
y3O8C5CObmBmJvcnLofelBi3yCe11xtEqDpUJrWvsnNrr4q9lT8cBXj74XcB3+kkmmw9/d35JHwN
OXPT3eN6A18CbIunf9ByUkdTgkQ+p9ZqQbQkmhRDUtrNv6yg0h/LBLj0GG3jM/+yk6nfiGJoI1/L
Oe7DD58eJeDxYvuZsYw1uFom+1cj64Uy7TLiDlVupOSl1UWGOhSSqg21o3jnSALEYhgp3ZGeR6rX
WpDXws+jJZWgZbKoaoh3wv/Nfgz58Y7VgQGGJmu29Xvh60blBUsHV6YNRZ5mgLLPfcC44yB9Q9bC
ol3btL+2LZbStmtGpSjngyZ9zTsOE2dErA9nIyYnTknu9zqNAE0RdVVIB4tlkL2SS0jrl/qoPod1
58KDcOVKlUQa1Ucv3vKkWUMJdwBFJyvpu/vvjP7nDgs1c4iyD1A9Cpn9S8LNSkR1A1XmAY9CbiZR
UnEXJ8njmkt70NCPdgW+lAt0L316zd08vJoMbCDbpauJ542h7koSMjNBTRJYD8LrfSfkZkIpT3zo
g0S41+QlY0YNa/SpKSb30uepzqHmzRGBBEQIfPCQX8t7G66e3McDiFtAcd5uF2FucU985aTvNi0Z
CqtT89aZ6v6EqU5UrmC5rkYHjyeQ5yffsVNFxgnls3iFqkw+i5uFXWA5AyWWmS9FWs0ZtaPn76pj
cgRuhMaV3RTtiB0elp4PXKPju1mi8rgGdlxG6hpTQVlxT64nLtT7A6FzLVSR/t2KXvfBP7Kza0C2
orxpTd77B7vH6EYcg3Au/IAuJBwlaxUfqOTrArioM/7wifxJ262rtJInH8WA5n6mRl2eHJIJHyNy
LRJBcFjoMB6sf7xAFLhQ9+NDiv5K7H68WkAyM1U6F2l1jkFNGtmMok66HuO3x+j23dzdMVlI6awg
E+2xegaIT0iADinSYqY3995q86b+tOk5zMR8OfKEMxvaxuUl5/M2bfIK/SM9D6SLUUXk8NzYj+jy
dOjAFTBwaG6V2/dwiQ0f7Ky27rtftcU7ig9JoCAmxbom9kU/64H47KMonudPwbDmS5Wor9G/uzs5
c0rxrGjRJB7Xt05j6ytXMNkfWw3EjT6QToOqL6ctKc4pRUfdjPc1JCt+TKV2jsGJC6M7CjCNvNmt
L8kpLlxp0h5umOlUiQFiX4mo2m8NDPvcLVE8LMq7KbCRL6ybTNEYw4zpsk407KpPIlZNgL/SIBL2
ULFyQ5Z6yacCZMQCZ04gUsvQFzQjxo6R8WE6teCxWtn6eXFhY+np56qBLb40ceHa9O/VSfdCWjE5
a2ZzTL4Ap7FxCrWv8kLNafjj1Pg6VJjiAEaLXdnkESnZTGabrp/j3yJPX9P9vCJtYHsBAyPjxFCh
qW4r/wPlpjalNBIdA8sTC5P7PeV3BmKsqS6XoNj3eGHcLtVlaSld90uuoG1woUcMJJ6G8llqiUHt
JNROju60hYulPeq9g1VUzzmDc4pC9G69tWpPoAteArzDoH8KJR2KFI30LQM7H8gY24UKc5hopBX0
ipMPOhvc9JGFvyR7VxEYI4ROm0Cb8M6J7aQOLQizF8OF0o1iEJ0i36pK8C7hW13fmB3AUvzn+0z0
9weAvnLn3Hv1Yvmx+BF85gTunlhY0el6WNrBhQ3Q/gosH2QnCMk4OePSG/OLNsJE/y3Se9JDlDRc
UBDpMFs1uqhxZkja1X9t9DIa5iNw3GNCGL6+3o6PqjIzIDseJzL7YsOM7XOgfcT6FYUWiDLykP1j
03KgrZuMR8ud4mKqUalA157oacopBkmTBAkuYyhkITGC/mUgGSyfeHCAZcIAgQFlQqAE4arz9WZU
Yjmt8bE/CkuWHiWfEjViJfy4d++W7A/3N4PhuShS8TMwy+hwC5ij87RRUHrqiiNRhtUFldwslgqu
qSs0ykBtwt/6t30b1XVQX7F2naueDurpCqLyzX4WDZCZ21MbcF7CswNx+UwuFqfRoHo34a8gTDxx
3LhFBzjFfq8jJt6iJEZH3y/vPTXeW6wwQ7Xck59s4GM1svocTmmSCgxITxRudV2LMNBW0TTE2W/i
Lcs44RYrwxT03xgSNoJhvdGNS8YF8ArpGLfFVcoF0Of52hymUgcbMhWJ6ohQBEjo9P+6cVCwNYCL
r35HHx8eC4fKSM+CK8GoIr3RdG2D6SqhR3WM9r6ygYR/71/1VbTywtttokeTzGKqEy/XidwohnyK
zg+mHX8N4b8+JTW4rvfL5aJ/VT9I+eB+7kj2N7A796WSr6UbJYH1Xw/tidgbfqN/oCog5GgXBaeN
DkUdxWYpXb7MAjgooKheNWl5jODo6kCjpXV6ZKTmaKbKcgW5+iTlc+8kNWzvmvGJ7u1Qhrr10PmG
yheKHczxEdml4GyzKmie0VOLLgSmow01jjCIJCPTvWzuXCY0ElHnipKSkO0pCa1npGn1tterUb79
WNh8ZXLtIv0JLmGKl+XUv0OgpK/iAGfCJQ4tqL4mCmOlsw8NzZJMOGgM3MZeRUx9FZ1MZGPIrt6I
rObhyj19iK3nGAb3lOEsm942lbcsf0j8yBorNVizbTX0elerZ0WI+jqdnOfLvV8eZJmHfhFoDfbk
pJkpUaPJPPUcTRVGUlLsn2vgvcPMldnEi/RFOVJgLkhC4BXww5G2Vrh7WOWlIm8qzwo8z+Au0qlr
12Gy5gLFQ8YR5cuzWMthSPYNxedUWfaFI9plYm9p9SR369iKE6V43HIUD3tcEV6hGWK0kLfgnYMj
5Bf9PfQgrqgh9jxJKYTVBaN/T1osx6zUzaaLz076EoyFTlVjQDER2dWLEJ+S7OBZfHhUXe32JYqu
y3Kxw2B6LM/Pz4u1V7FaUQRw+Pn8YvbmJvtmis1hiayNhmRk6OBxYZMOe52am49OHIefyTGCra9m
mLXH6wrLw+mW/IOtIqK1PS/e4i5o8CDME6d0s5bkkLV42oSZ6+vMBO0Q63wpK3pdDFG8ORTo6Seh
WluQJCUgqmPjc7qfFvHoDL9S/0vLwz5GXMk9v7yqHJ6P9bJt+G8oAt1dHwSafHGcOly1e7spHmrE
Vmz1TFjhTJkubUV8FJhHqS9FkCsW0pD3aBf4lX5B9TI8iUOuaAWXtkvEVRdxZvbZFxeCxx0y3cNz
Py8hguqX6VDU8G98PVdtJcOVPM5PLeLvFM4VIn9ntwLcjmYXItmH9x5JLokKmbrqgq0zMQU4GEBu
WgrBtBvizUzrVkzmrk9Fe3WcR/LT0UeEsVgPuW6OxtZTFPTczHkin8ZWi2D3YRLJ5SGA5A7v6/HJ
5Imv8fa+ZO/fjfuDSSMb+P+1U6upgXjdMtVEPOCSUrv6pY86y3CwClAVjeiY/NfTIQXknTBCQ5qL
NjdKcsQq/u7RNF9RjHaNN56vhM5U5RYEoE19zzoAsqOdPEcHZg/D0+znRBdEjz0w3435fcKiXolK
t88EEMStIJdpsn4vGeqTQ3+YPyeW0lGOyfhqqOGXNQIJQs9W+c2RYiyWlGvoYIMpT09tRACingWs
4xzTdQvCu4obiAD8rmv7rcSh9zkl9Z99qn+iYCniLUGv6eRj/+lg7MGognBjWRibaZOnHZuMa1td
cwYR+YOTZ7JGZIE2BTZB8RiJ9+xC8Gz76kPkCFgNW9GzQ2CyIn/1WOOU6kNwo73vSAesLxozBnRj
gnLhjBWc7urPzRJXczh6tEq3Owp2I7jawpzeSmDrLb4qrfmpL9TdkDdIMoRBumm4yScpIiJ8H8hs
WZYcND5MclN9oBNlvdEtbLQhl+LbJnvqBaoCqBVfFvBZ8mrvgAUe4o4xcJNqQWfARl8TG226RH0b
4c3dzm0DO0a1Ndz+dMdhbyHQW9w1RN+QGCgWh5HecreSr7WiAvGFu68muGASq4QN4aihtbFVns5B
japJMdyRsnGFF+3Yi2LBph8LFcot1NXqTj2EaPK2eFAzGSaeW8i9570HQj/ThSa3eNmk0XZBvCtH
rrzAzi9QZK2jLfA9T6OmJgWw3sbvMx7tPUO3EGY4xbcZpn1gOq3hTp0hS+15529I5E6dfMMCug4y
UkxAfWaZ7/yKGDCv/SW7hhOYKn7thDqmWflb0yFmSv62foFYT+Xwx8TsCcI9zJnTA78MiHtg2iZ1
s0EmSbgFdX2uIKnI+RzJ+1lpc45gTGyQTKl/OHPAkVNstaYHQKqGdrA+GD/Wh+zSXmyNOiGnmSbi
uH1/+0qgMu0fucz/p5qbeKZ82bstq1/4+dSnbf03P4QGqn13FGEz7Sm+m75fDhEY5px05wC0W0GX
ysyb+un1S9YF7A0Tj76OVerEM9igSBbFmkrRIABx0PCasaL3WRLKhevCzQrkUNtkmgmMKJnna+2E
md976CcSeMn8fLDG90dzFZsYT9FhaFgjHxiAkVK/73oBUEIwLRCUu23FCmLfGBmCHIe9ssk89JNu
CHJIF0L2ZIL+WrV8DFDitzUXpqKXPDl1A6qvAr4O0hmkpVfZudESZHNjkTdACy6i6jgEEhZowdnf
LQjYs8DNxydG2bJWQuFgYcLYWpSnmf6WkFVp5Dl4ZxXuUUCFQNYBHWfTTJRD/1ouwDR2FPZEJaND
NlDfhVHLnkqWQ7kfJWhijmwOAJqRdB+8/8PehxBEAgtg2k2+Z6NB7bN8poiwpW8G8LNsO7EHms0E
HuB/cncd4AiLLBc/xQ4HHmozeYn85cGliboHLDrYRwAB2sbrcREugJdwvRs/ut9qQVpLQC/S0FfS
bHxYcRScb3Nv97KsKv9kQGzh5xmpDohfIxzt2wrvmnw8NyJPneT6nvFmuvtQNkrqw0JC1Q6Q0Lrm
4QZEgkll9NlQxatI5o+XeOn6Ax6Xrk7Ve8HdSsXZ+q/kLfaCiwCrlTg4RGGV/tO2/Th2q84YBfPY
5sDvly/qaA2PH5EiT/cnsxH92tbC3VNTZprWHJ/2XSGpf9pEJpowLqfOmkTyjI/LJnoaGGwbN6jP
DbNwg3JUjGGuXa1A4hb6A1qZ7vRLkdmdFM+Zno8eySXErOnM/RE9uoyRBfGIUr0voAudhSNxVteV
7WeURSqCecJlwD1y341dZmw6sT3/vYOWGw2jT+bACScyIszLVsLA4RADdc660k0Xl3S50I7bYYNc
g1Na7zgFoxIv6YuQw3xX+9Frr30ubzC5gPxavsZsTaJ+3Eh4V1EpBmN3r4Y7RjGx5vx79zqiM+J3
KLxQhpKO74OJL6gnxvL2Y18uCCld1LNwYHcsMf/XdHGoNW2f+kVlyJAaNThbV0hmtX/d+Tu9A1ZW
viP2ALdKBwHly0Gjcc0jmthrzn8MxOIjkkO+VRw/r1sWJ2md7MkwKX2WIC0re7+Tx2MMHKz3OVOj
SLIquH6k4oXhfGwBlycajbOByy24oE4poUoAQ4FZjbTzeuuO5A5fN4Zc0w+jU9iFebBZQrFIYkEV
xulaT165gQQOqynJ3+kzVwhcF8xcB9aHmKf/AvJjfeS2OKbU/bQ0r2r0yKa2zjLDK2cLdUTQREsN
/5uVQljD6B5uPuTYnB7rZRWxGEKiVGGlhcyICn7EvHjb0pO3dUh9e6/9bwn72NwurttncB03Tvyl
1kkqyvadhgR1gkocOn4BM6VRVOrz1aUmZAySx+55L+K6YAsYZ/y7RJqddUhYetwIEgF9nebY+qXH
8o2hC/xZil89jIfEkXntHM2W9zA3/OBbj5rW8rPpG0G88TGiZTIS+7DcCPAjwFFOr9iVtitHd+1K
wegS/XcJeMF6erddHtCAWyvZtrIp/I1zQBoSsXhQVHeL2/pDxBAxlXSuovzeG50QlkFhR7Cw/iYE
WmSH81qqpfNJg0GA5USo/uZfK2n6q1C/hGz8HpwovnZ87NoinxA9od/LRbu/Q4tv7JcsXlcECCKD
3byf2O+kV/eailKWFpj7TyHylRVEVsVb3hHFjowxqJurcEWr9jH2fN/ew4HTiF5HPmNP5skmJ9sY
+/ojNZTAgcQBICSR90imuKK3Mxr0dLOvrlw5Onx4mWnaCUmu9zbA/7nTM8sj9dG0AyPJdxuOlxeM
mSNimfJIdLzNAuRIxZUriCooYf0zpZvSep0Efz5ptCIQxjNQ4dnRVRMW7sDyqchO+hBV8Xc4c1Gq
odEJCn13odYxpmEZJoACvE6J2WCMheyH3S2WOcDeJxXUQIiIEDntlCDXhJXdqzpS97IXcLOdVoVG
x+jjRWwrWbkhZiss/49CT5xCpeX41eaRmr6P8ED9jYXp1GFF9Q30orOeZ05T4ZIRGuZXbAkZu2Dm
n6ci5WD0h1V0hKdhi9nMC1amR1+/bl5a+P5qTakBsj2UT7Ur9L6+0rhJhP1kt7Dag74UjhrY/jqU
dOpoW3TvkxHnVfN+mOn1F52mNnWfBp6w2/qD7RPxjujvq299cVUgbzsfohE9NkKIjIniq3KfoEze
j7jhjcKTU5U8ob0g9R2ANweOoSfM5XWejYm3znWuBoQt947aBOZ9rUjhyeLMuuldhnydTXNUygHe
xtEzTMr7S+iTtoKgMCw6U6sKTSvfnt+MRwe/vzFFSVVnFptDuczIai37e8w5lNFfMyDODdVGaC3W
A2lQZvDpZuF8xO/Gm3d47Ipb25iC7ug0jYd9gH18ZNA40Uf/sxHfldbjNvJd5cdCff2eEewR56TY
JWPLvHly6MiMgicqwyzqAlv8aorokn9885FpjQJHdrF1j68KiBIP8EiBV/DQpL/tlsgCEuQ70JXA
MG/11MCzZp4hZu16juRrsibUHHd6Y7dr9k88YWRGsOoo+kkEZjLgTi57CwKSZ8XCi+Lny0M/7+66
Px4Ydfjxb03Oizjxls6pU3B+OnJG4eCEicP31EkioRIWHqmouPwstPPVe6elAgCa5tD2hk//SzQs
eEtIdrzoxGAfgwwu7ssr8o5QTB67yfIDGf7l+jXTX4zEd58V8vcd4+NYigQDtxqAXvyarBhopEd+
v4sEe7TNsN1oYXrI1miqm5CrF6bd1oQLwToElUxPafcDAPne+Gpel5KZHDfYUXFlNmLJnURd5rME
cE9q9dyRddYVtX4QJNAM3CyguDEVim1TuIq9+VdUIjZgDfvwy2lB/Pyr/7TmLrYVdFoQwjXxp4Mb
6n0SqTkPzSk6cnBgt83ZQ8gk0e0fK+Qdt1udcZWKMkb/8b1jBhXZVPPggwjn6ZEorIpN2GfVXGdk
GuRN5ODfckapH3HM0NuuU+z23CSwZTOXPailr4HNn2boazPcdhFFGc9WFLwXwFU2EpXtZr0IcbtC
+n2S7iX2PNkaVfS5aikKyBlV3QRPqsGq3NEyZgNodZVMjGcScEcCU0x1stUbx2v0jEz+AVeRkJLF
NxquQSDsny8CgMhZqYELHMiI5gwdSpEfWTN2z9mk2rxRiURfAajh/QOMp8G6JSnZDW6hhS0qd2S0
vt7ujoOoosnd2Lp7Ikbh7YsdfHMNjjrSc8g8eYlt5t4k0tHln4DKAX8deA4FaxCcYo11eNZWLnkx
gXKZ+xUkp5pJHOjKQX62Lpl9spZpcEK780BxshIhofyuRJ7kvhVaPkuhgN3FtUqE1PK8wX+OyMmH
BdN49P9K/kvp0zPNG3tXYifBe09htVXTdUQIT3w2c6ynGFcgPO1UZdbotpv10vhiO2eMEHoFS98C
8WPa1OCtRzUXVqsH+bXHrM/yFxFyhWK5Sa/hGnjR3AnuRzBUPbw1u25rFhiIokm+G2ol3TftqDSS
mH1VTg1ZZCZa3kD8QTcyXcUBJ9Jv6aTvUzuUDOUjzRywpOzXsTkrnOgFmq97aRxrAKGVqQxvxRcf
C2nrzSGqUTYQVIWRQnXBHJ3CDlbMgT9kshebZ3pGeuIZZOkKN453qrFHqs66pCDOjyKnz4ItduH1
V0k/E4/XWMXBMC4MpHBxFXJRmfu+vGXnOMT4f0KgXuo/sLv1REUOumXRVOpKTDK0oBsodhNKhLQU
m1CmNKsslf8pLpXTtA+4SyPO0mmMApuSO1J+rd+8SRI/fXTg0Zpp8I3GxPV3QUQ4H18SC5LtT9Uj
XpGaeKHD4km+Q1nj+vz8u059r0rwnFRa1OurzfHryREqV8BfFk1VyWSgg4X2v51wOpYTD19Pg5WU
UW/tdp/sJ81LmjL4p9bmIQ2PhVGLvuSQWh55gPH7eTDeJP7h/I4iU/+6u6M0tyF6ZEYM0pI9lMBU
gNgr7zzZd6CCQnkqxjR8FtAi01/MBqAUGoOrdc7IhnuOtZrUS5SBY3RkFA6mj4/YoQoQ3xVDDYR4
3YkzxehuaHT395UWTg5rq6ZeRIkB9WtWNC5wYPjXHVRTUuvGRQO+buZMCmjMulXGcASgyiemIeyv
g6rkgk1GPzRyvLfxborxhngyVgersyVkaNc8BmZe1gz+PQbZp8fNEEXXpNZ6rn1YW1hYuSrzpso/
jwuRgyaSsFs0PorUdfieqhawaUKQyTGQH5roFCJtldkIO+AgPL1LNF097S8LAJTYKVbKzdJCPIZO
BGsMTjuYh8nvMZHT9ztC/9vClLtxt9TGXVtDncLlByjdD8THObCidGOl0FuX4ABQvQaNYZI5mOXl
x+/DoGjPMhUKtxxjkw/jIGnYOlMjCvNhsZMMJMFNS91Zz50WmSZrNW7L8snofdqH7biS40BSLPY7
4zDvAfRO8ewTFEBkvwK7YnL4Wq9jZmO4HUoxdz13StsaZssJrdVOh+FZw6f/0nYorTh6RHNT9BKY
kaT4tKYrIGd5PpHaTRo+NUNna4rEz0aEWPtnSViCJ1WT6IEXxyocm61UnhFULqUzZegKfaZvLtaX
SZdJqEdjIcX7TcC6W2ahnNvbpWFzK4v14GZ4wOyLnb6pABCfRI/2BfG5eyYcVX+P9jYBK1ARasWn
HW1dnrjmnP51UhpSrojVKwrv9iC8j/e9HZOW9/mTm4Ry4enA6SbQ1B+l54UZuhwvYf+XlMEI3X6H
raiaebcvbvBUziJJjYB2O4Vo/2FZ7nXzs8YfJO+cT+CvGNs9EngKBFziTeICnpxDEJVT9FsOc7Oe
1P1s34aTKkRVAu5ZexFKaeJy3I2sq7rV4KWzOqmQ8PjY/kaDu4+jEA081qaJqOJdRKz7N1KaSC+M
KAN0yVXPhlf0jchKXnFXBkXJ3wnnoIcpSxNXyRvWJJvsWLl5REamcuF0yfZEGyQV4wa/yNby0gXK
yJ6UELw9o/NA/6t1srvuevd2mE0CIQ35vwxT+zLT8w5VJaIlJeoA2cUQSehLbQ6iau2my6k6b7Qz
BcgK/CMtiNnfIQCmF7x7Ui6Pjm708G8839BIXQvSgtaPaRFskClrwXjfegwRpMMJ45vdO15Ckh55
ZS3U/cKsxyPszGPVTdG8Fw9dyn6whAadKV954SBAm7cN9lLZCR1izpVIQCCHBqjKA25St40yZvXZ
7Fh5yFHI3OtJjXrKR3TBkNzI8Ybdqqe48hni4+TTLOkydVBEfzbQyHDb49agS7cMNCAuAHzJIH8o
UzQWQqy4426m4AbzN/ZvmbLLTjmups/SzgyTfO6y5vI3yi4gBXX0NDMh3RITrTmxla1d1jjoGcFg
8yh56i3feLsF6o0DhfCl3c03IQS6MA3PBkfeg4aQfF4dtE+kV2xCuMjibYQr45x+Czzxdw4BHeRS
fqj+hc/2WR+O+ttdxkdtR3mD8ffeKqt3jolNPv51vVWLhBu2Lzz3SP5rz71lH1KIhq9wbTrrSt4E
aEnxc/GWlFLIQ/xBYXKvy2khbiOeOi0biQ5/7sJ/2b/Sj/FfcKgHmy8vT3kcQCWmerFSJKkLXN1l
WjTh6tVkzA4SwOzbeszYNco3hnBtDXNXTfJSYYBsv3f2aYnPZwx+cBgfNSa5abbcdjJqwlSwJpT2
3UZPX4fGPn3nSoC0z4n6ISD4QRniV3in/RTUYZGHqKNitRqVuZA9pIpaibBu6WS4jc0FUk1VBZjI
QNc3jqWBHFNc8muC3WciPqaEUlomb4E8VZdQPp19nE8Q9ZFchwdd5//zoAGGe1CVgijxR4gIq/sK
rKaJYZY6/Zag7lDCmBIesrk4KD/QdTmVgIS1/Jrma3hATcdwd2Xm0If2TtlXDND3lbnyInJQcKuv
QJfHvXfhGAyvVEwJBkWxyspoW31g8yxm0PzIKwSYmlHzEUiFgj1moASHFDN49E113uILfEzqyLyb
Uu5CbR0F1OnOBKzhC0o+hBksFiGHeVEKcX9jxYSEn/H09a73OTG+C4pnSzEJwSN7BVg5h6uzmU99
8ichPHaPD4ohCMLNvyzp6N0IAcYwgnLllPzKo/V1aflDKJLNQs+alp17dOSJm1OGtxti+7GCxLm0
Jv9lW8Q/qHmafrS1CnDX1PLctjKzYAhBMPQZi/BZJvzwE4YFrMKTdPhYJl66Wm3/2L70gzWUPQtA
Rcx5SepnFEdj4tvkEceq5HhhHkmZwJZpnOCIEyGSL1MzjpcNkolANr6QtpnMy6K6XZslrMhr2WJc
bcGi5ZR96Ir3ZBVQ35K008bylLA4o4ftv4zyi7eW453cKhN5MrEKUtE5jDmzrkvo+Gw8eCjEziBQ
heDyY+6HMeKVezBDLgQOUPLSLvOhxGb736wX39EcMjTj2xUYInw7YILj6epDjYCnC2bTdbOPCoUb
lu+peAFjKZuBTGYrDZYnhNvBMjLm7nA6OxOQQAWnRo0slufxwa9PSpEIqcOpAlPEbVy4EIxb+gxO
fw6QqGJ9BmYIyECtc+wFQw/Zue2fDL+s1dkOThFkYIl3zyba1B0yicdZjVp4e4Paf8z2IrB0vZxC
/V937B32aV0xAL34RBSBcxeNvzxjaYqLW5PudF+9TlgBOfzlNAC9JQgA4wDFYfI5PtAoEvtQQ91M
8YTtSKnuG0YDi0lSOaPQtM1jaLmOtEmC0yz6iKn4lxh4OoWCULfZ8+oXVXyLB3L1m394KakwF6uD
nTXPEmiaR4UpkRwEox1UZCqFTLh6/H7wGrxuHXUnDFGDmX9nHZGCgpHK+Zeo37gnmn/a40FI28o+
O6KLrlRT62i48ycEWKZfW2X9Vsb0XKJNYUTKr81hNAJ5Nw3Z9yKcA1uZa7c9ckNP2PA4OyepcSNr
mkQ007z3aGgxWX9A3QpJZlbjki/XaQU9CvMdJuvjfQPzcBvF8nOvX8NqpLr5v8tPugAjhZ25ifN8
EvM9c4mtmkKcEm5o7M5AzZFiaolDLLcHiuyfFtAnFn+oJocY5mtcCx5ay3GnME4dJNCA5felvvHz
eqTiEKmGRY8WJSLYmw2jjm2qJNsCVmoBYifaFp1VkW+ugasS4S9DqoVrgPPySlAS9gfFV/1eAh51
RWSp0/bb2asve2lHOzcLK4Ux1ShYN4ysC+E0tiR4eN23LA+LxR/02FpdaTpSf5w+pH9cf0Wwho0l
rH3RUiURhM35lyXHPuCwPg0Xqhff9EFybB/o16myfVjm5NtpoP8LFzb0gReCPrbfTMOf9JkkVvrD
/gSWMAt6I6yWwDjWcOjQYcBiEdrK52GWnKJ0OwbGdgl6jJ6ZMO4WWN3UDokZtePDjX1b2XLHgIyU
S6AfkwOsLuS/dHjeJQZkdq+skjeidbnEpw+nyLlFZA3trFkYkp8Du87H1oYGNtv8ZgpqfeJYd2gB
kEmYxKHQY1tYSYgVe+UGTyY9GD+8s0TP/7Zz1Zk3gRMEkbryOcwd3hvDEScrxvhpOEhKKGE/5rRN
jgNEqljA3EPrdZ+YyhH2cOaKlpdVmaDizQmdJGjKnawaU2JM1upJ9PkVfSqoJXeFO27XwcDEQUJH
ppBdYcmCU4/rKecuRv2yt+58gcy5UTuCuJbDef+IcxQ5/bETxb0TvgvNwfi4Vs45TOe1OvZOcpYr
uBixNkaum26xANIYpeOklo2CuEwqJsl+15gJmAKEyMVTy0OMHHt0KEXURKBxg88AQrd1xBs/UY/0
Rm5gkCvXhpVDIh0LUpwD9DglBoNu/VrtoOQuBIX9084GsVHtMH0ZQhPddXMex91QCDu5QhVBtsKA
5jpUB7MmhMtCx/kQ+1yq3qOnWJIydvz5OYo8v6wJpbksricSHbaT0zr3Of+ABhPUO1cJwFaWXpJ8
6vsRRcuVzkQpmLmOZ6+R8pAI4ADUfMDK5mPwP7+RwaXiMn9F3z3qr8BYbteQKDz/gjxCYf1cKvVG
gN5sjw/pTNELsWMgrvqcL3+9TWfhe1hBWC/mctR8gGznVB6Csa9kEzh8rA66T+gh0C9bW54M37Un
JOkKPG0Vx/VVmFpVAlOfCYtF6TbQ3YWSZhfJLJMNvTmhFq8wW6OT6Eg7oMG3CEnSasxt8Z7LMmgU
dIEmsrHH2b3rIrzR9RFf4OK1cQHCT7POOB9W1//uR9QYbtP92e8T5YnaIOS7QcD7hoaKABRtdSuh
mOYSaki/pYG95LnOOID8+OaRHHaO7rd6wzez6HmUJ3CxP3owfdlgVpaG4re7Tn8+76+DhqZTBhLc
YGVEMVl5QOQ0asR89SnWRkz4S5iYJq0Y7rfQaLnBmNjrEL6O0J2N19SC1GPbDNl8PDjv8eBM75Ak
41mUGytG4mAixL4Udjw7TeXT7gRyfR+xFPAPGcreo9QZDlwYl3UKAQOFiHPhGAlOjXcwMU+wjAQ9
hRb+NTz83lQb/5w4J3/c5sCJMz4wuQSnd+2wJZ03Rh5z8jgDWxN5sLwGudEmzdTZz66fQOUfBvP4
ugnm33ajSLH8C5KO6FE1shSrmRzFfmjcTDzwTJDbGmGCblWVtgnr75bpHj+Z3c2mee4VIYTQDx+R
vyl+DuvBZFLj93HIoBa53R19rnPh3mTIURcJFG0tY2O/Zd/g6xrtgNQg1jQz8iF0nlglAFBzBDa8
CzAcPHqw6vyUUhF0rDZTfoUDJh/BVjdKJpTrkeW/tdG+py4F5eOKm8Pt7VkEoQOb2rv0z4miKRkZ
6gIX4aUVnm9dyxYe36Mhv61AdPMZemMq0F/E41aLdnTmGgt24PefHQ+41pUlsMHwjHpT5li3mhpD
X2VQJTTK8iRI12tmy64H33f8XBkP+kyUCFvUTTBoLAn11kFhCXsZNp6Nf5pPXkadvQ8IFl0z2aTp
1LsDh34kt24FeSYcPyYhXkF+ngdi+0MdBJEZaR7mz9jtFo2FSK8Ld/XZVxvWl9pGixR/y81x1hYF
4U5RSp6SyuZTNPh7Eo+Lz4SpCEG4rQ2Tnj2TPh9HUyVmQgvdnZLqWfg/4lhN7gzMwf3cfczYzvQ4
4W9gGhVRcckCXVizR9ZU5/EWhI17DuRRfClmT56oVwVVqPpWB3zmlHgJCocnwLIKAkxfb+bUSBo8
Csi/V1buxxoiNmhGMvOFtDzl9A/6oC66YInTBF5yMDAl5dP3BSnm0sB7q5UQFrlN1ymrzBHW7JLt
zyKRNg1n7pUnzaCeSD+vnQLpXHvtTugQfYeulCc88M5tFocxLQtLD1CXDbx8OJ+MuusxT1t6s2qe
If6dQXxh3xkdAI5UID59JL96y8tyYqwbor5a605s2vaGa57vKTuZXP/Kmt9xv54hHrmEkj9glw2F
wa5DIz8kVPvRv0yChMh5JxZM0O0X7nwy6fH9KZzwh6vqQerj66Bre2eF1jJoAIAN6AW22hj5RKal
Dhv2wSeF5VhgZdl0dinKWgZfNPXHhybKI8t5HbX6KbRY3onBOVSDw6U10NDvhvG+NOSxjq1S8jAJ
mEfjBBs3dkhzLwv1YulQ7rH6Xq50su686gexrKgUOe7Bn9J/7pw6uXWR+UAxRN2CTjXTrKUg2UKC
9f89+8VTtqZ5FUWrlp2mNern8dd4yI6fK5t7y3Aob3VdQiWNh5axcW1tAfTSk4ZxlOS1Mb/WuXb5
4tI5n/QtAJrT+jaDTe5GpuCSh3e+lP1+GSQS7fMh9wKoOHOVNLBCT89SeJ1O89SpUiQIMmauHuDy
JGXXRM8fHhgEa3yoj/wWEN1c0e6zgUMzWoUgJVkdpDb06apU5geRpyDpo/irZMFFtL0XHOGQXTD/
XgIec4L/cGOb7G0K8zirDFsgokeRT5SQPxhjcghuLuSH9K+bBRR3Nb588oPOAINswksNu5ZJ8xrA
a6I7GriN0bhkEf7tto+CIF0QEnWln/f/8XxcYnxjgbXr1er9RFhM/A+v8noccvSXdkWVlQw7hxGB
Q9tcrvWNfRkqhCwmV1v2CF8IN5wJWTrOtbWXd9cP1nYk0Qv0XPZViscGZ49z1mBKaMevBuXVacjf
Us3jDD2tpg1osecTXR4Dp/5r4y8SvRR2+yvWIEgCM9hyrZslho7/JudeOMpDASRqTCAQHDw87Sd4
otHTbMr+kF4rTOEj/GFoKBTLhP3SphnL7S7cvSzKJ2YllCLdYXt/3ekDmbh2Vekk/ivQxuvGbKSW
NLDtSJZ6X4MFSBnDzsw201xv2ENI6aaQC6cSl/YCf+0ni4kUyuNvhMHGHeQcQ2GseJ+oNod4TQpv
gtgqsYyp0ULEe2DlOGgpjj5O22/JNo+xtEnR4InxYHxJYVKfTjYnAKinyQFDw6hDumO0zf5BswOT
Trx1C3Mix5i1iHjKbkSjqTnXfo53E63fZCUQgaj5FbS8ceHNtqDu+I7jgVHuam46kAMjQeg7LF1v
VBgenng+5KmptXAMGUz6Wq/KdEpPkICNyHuX/LJuckA7C86bBvotfxHBzv/SVoKtMwGdZE6jGAzd
tgpZp+UsTSlEoiO7LHwswH20QUGa6gKbpZzbGRL819VdpYFkNQulVQD/okFJZqQix9+/XLioYrmM
0tNP6Khcgyfe0vbDARY3KZsL4LTfa74/2od+TGLtgYYHPd/Fsu4KHY876uzFO7DuX8UTQ+Da+ipM
7MAhf/HTyg74hlgKkjEJjTb817S2usd4UCPq0dDmufxN/Dd1iAEDkUhlnWLfoDzocPaKrXQtnqQr
HC2rPVBCjyn5QbwdugKlcsBviv+R0/5X60QnLM5ZJ15vI4AQCl3t9kRLOQtsB67/gfxlIwbbNQ80
gLzCb25r2y7qOYTfpoqSJu1QihUim5qYu0zXm9kH+SOYFfpOreAUD2VgIvtyRR3TjrOpluWeg8cE
6W0M0iCvFXBQWCN8YHTZ28AF7u7MJwnuDivd9uU+eZWOGGYSolK8RahWQzpr8wUFZJ11qVUZeNs8
Icf297j6sEpDkoxUOQ5PneH5ULtn/4VSL2UJYm/jxa56qI3OEaUQZVJ0mr2MwqphX3lLQaFItrCX
kExheu7pHMi1fWkSMYoU96Rc4HizHn6PygRsZYo/1uKtRYDEsQsHecyjaOOOiACHI2wNdb2CiGfo
9XQYS7x8/RenLNOxli/lgNedhFk+X7NYHT6TDovTy6zuAiaaIplhC9IWmmijDTV7fos13E8dcqiW
JqyyRHQj7txhBo4zLocfjlLBwRmMSqUOzSUItwwHhqyCYQKi/12tnbWFphQXDlGYapyOKStF+ta7
tQr34kIYR9baJ2BwZG+EqDM9n162v+4EB1SDXh0xgdRZWWVfRiP+gnmSUvz+djghds+qfblga2ai
LiPeq8485xXkjQI9OzYjaEILw6Rb4o+tUEr3ruXPNBI2SYtGJ68jmy5MGmnbLgxFpSdtb9yK5Ww2
vdDBcojawHczGzKP6nGgBDhu6Tdn6t3lF8tWOLIS8Nul5E9cnJ6y8P+zdfPT/WGliIz/vuOjbq+T
quDBCXfOnWfO1cFnvrcjAUcdZ5xnyIrirPYak0Bk3r5miOzc+p231i1h0vg46p/h9bBElAInipOu
9mk4Wuth2895XDzu+goADGrPsyFEByFEPe84Cm1ss9mMvb12a/s/yO7qtbR1jyrn07+U+rCzIGtd
VfRUOCSFum8Be+qcJtjPyiudocdyMYjRkbsXvYKWwuTDj4sEe0qd69OMtW4MJm/zkl/jiOgxW4aU
Rir9vpasWOYc4jd6QFJZk7LgYBdcG3UNza2ZUJ7iE6w2T0MH1FnGjCWfjm1U5mKGD49FXyC0iH2W
KVarW2fPNjaCDIpUUxVU+wq+dM5hVLKKJss3+PI8qaCfMZek2Ep73M53YIYmt2bvvvDBw5cP+yzS
lYydXlbPXus6aepyyHe1tCtOnt4uPoza+dvTcrhhIAOVjHHgMgtUq5orUYiqHxITqEOgSGyc6Chj
HbTXy1cSzrJEArtgOfP5qVDCnBlnRY/CwrRqev91SBuKVHYDhdyA7g3gbNXmagZ4A81P0ebL1aZ4
UKDRxZ9gM+EIUh/3ndbQ2CFt/SSnK5FUP/M1fWc8ZuI5CNkgCdQhpeVyqvTZuCEzgUgs7zwP004V
sNHosBTzZ6WlYmBn7aHZ2W4sDo5wUy1yuqGujSG1LagOEuOezcaWw2U03zZM8aW71fx3SobLULTv
mVNtJth0xC0dSQIvCtaAPHjTH5q9+7He96blEkTQSvAUPrzWwa3RMwDoS6MtI172mE4r5V6XnNb7
+gdy9P48J/WrMTMRs5h0UiV4nAOk3UlT/grzHZXhx7fWGaYz6lG4vF/bWgtel5983Yxst39fXedK
4ZUL8S6PBlSBV3E36UvgE+4Ae+XBUNmKt1KXY3a4/Oaaj6EL7vmca5/gfJNoQ3qaWt8bg0/1WOg5
ajxVMH3AMyrm6X/ceX9DGkw/0EAIbTCya2kHIZU3/KSuwdLl6758hXvqqi1PVS/vDEsq6dQJ+lT0
meXf8ix2tNV6qAKgcBYrRBxhvO4n0a0QB+9t1xjLuZShzyCSy5QThvF7nVgyjEL0NWIvsTtiIke6
vNnVyuAmD9ucYi3QfKZo7CojNO3gkvqQoVlp+VmBhEVhw9VUt9G+2tw/r8ZcC0YagUw43ThQBKk4
/dStq9Cf5Efgqs+sk3Bg1ZoUCfzYfOR0j3M5b9VQVSd8k4gASfprrUJcqoveZlMHj/4uaX8Mq3Nw
MadYLdV6Zj/PV3AmahJCRMjqt3gdXh9R6rHmauGr93rN2MY+pIFL5jdhTyJdt5RCafPxskgY2VgP
vyDWQt7o9jgNJqz1Zq4zQjJf3OqJtZEIyMzbfwTRa2FjW4sV6oC4VZMwo0wuy+Suk+KPwfyCrUxs
FMKuzGqfMykCWWHLho9+CBxzj8Cuzpd6xO1IgV4AVKy+wStLPXDtn05WqvQMkklm0t0spXkIBXbk
xWOcZSQua4ieNI7DR9OiZLi8yNdiyvjEuYzfU5eBLzHXw86mwwzTDvMgR6e8eFFD6YR3mYaDtYzd
F32IoV0BQA39/7tz+f0uctpTjf1OuClPntkaWCcuY4FpQC6UVPmquo3xdv24k69Nncu8n6L/tmI8
phLTs5MJzcAd8x/hPwmqHBaeThAecbPsQPA6bzl2kyEC0RkJhgmmqr/oI542NbvtDIrOVj6JHkHK
bVTb/GdwMEm1PTWiurBQvJCGn/KijquWFn6Dya6An7i1gFXhXmVxX41mne7rLhR++mgHs+askOFN
mXfGERPtrfrQfYo5AGZq6mqV6a+TvVS1gvo+hoTg8KFmVVU2UkotC2x7ZlhEDcTgQC6pLQimaXrp
8fJ7XyP+pZKQv5JoKs1+6Y4Y5evZ3JT0ZYd2ZTYt/cK2AX76dTcBaM7aHt6kVdpChmEbSxzvICJb
LhsHH3a1J23p82BeaIGZiaBMm5vOMSW5i7gkVa4p14t8Gxt5BXPuGKrzCsVEqrO3Mt4RE+mM3F6t
RpZ49SSSjptVAFxVOoYP+c38mHrVFO/vsqNss7uBoFZtW2DM1d6pySuwXFQWV7FuMxSPYa2i3Ltq
QQ+d2LgKusT0SMq3k/mSUpGDPhauALrQ5GWUH7vmK0c3hvTtT6/HixvDuUNXT+SQXMAGNUko4Sjy
N0HCphm8UZMJvonCSYqIRVlIoWGS0M5n9UTUppvndKrNiVkiBqW60f+TZZo7xssYofTiZy3epcVS
P3R2teIOmTXSVy1Up7NGmLkrCZE/VkKGRiGJwWn4+ldXmyJ1qH3HWM1tmWuOxBk8xYWFFH57AbJN
jXd7nxCLNV0bEmtKRNmOoYbIUUrOz7SLOciNs9Vz7V9Tv2gjoeFKg6crBQD7pdxXnzeZGcw8htwr
VbSukE94LeOa6CdvFK6dj0GS0b7mDcn8PyCj5BNY8UX8hor0gXthiObslNiERckhWDgvalF7fd1D
SX1Bt73H7i53GKL7ehFYl/PnaVgBITdy6QXF+LzXO/A5qGT909V8mj+4jjyZxJLOSDqbvEP+lwo8
ayMKamXAF43UIhmvXG9/KHN0eH6FujJs5TsXW2vNATTnYDJAuwI40oVq/IhXlvrxQCLEAnu+B3sq
UnVjRk7zQynAzCO3xaRrLhmtMETMCTbO0tQQkvHdXkEEP5UVxUySuSGw8khEcs4LZolJ3wsKeNYI
yNy2s1SYS98Y/pYdvfq3G0ZotnfFXqcPS1YQsCXbK604ZppBnMu5h7v7r58QQ0jLg0tytkLnHkZE
A89u+7YAQmqgEQsHjMt8qimlf3P6ujomVjkpVKFffLKtk9mGe0AtXR2aI51OufqT5Yn2XEvk+J6p
/PnDAb1985qlZjah1iNtDZQJmR0K7fkRjL9Zl02dfzKJSnJe7ATlnGXlqDo4yp4LOCwwHKXMugVA
BeBKTfiQbXWsAactVEqPmRk/zX7Fm1umvBcKJcK5SFewShrYx9AREQWMh0cGPYg4zz+M8CoORQGV
FCA+emKj0jUcv0+UZP1BrcMFRwO4AB8V0FydabS9nMpJl23Sqjd2aGfwnoAwfiI1ouk/zVdZUAcA
u2A94004NC+EVDwzx4hdz7e8UDNEhAKyBdDGiOk3xeuRhcXCwJrFJn42wufTYG4YTEKsIH71QBNF
atrsbpB51bq0bJgonl551AN7qPlPBeQIgPSjcNGtS88Gw70U63HDRf0P2P082lC6ZOdFEvXz9zd/
2o2H8NO4Ov9rorU7m8XNdJFdCbf9wd+A0q7om5vbkycTvO60vdFDPF8iIxftklYbfcqlPr5eZ1rD
vpitOGWYUyCqbgugQ/JlKJ5oDfUE2dbofFdRB0o9sMIZ+1P0qgPbRmAAb9onzxNK0HVA5vvqrqNC
rsDQbesPBhytWaokW0WLGApcHz3oexiJxzC1z1rEJjh8yFGVQqfnvztrWK6DC8klG5QZLITERk30
QahvlllK8Vg697QMTforc+86kahTX8+v0gTks4ZQrOUh1FIXxHA2/WXf0KYn2HpiXUINeGNhQYzU
g86j4StwANYXJ5J8CpF2xjk0sb6tuVnWSd4E32r0EvDXsC9SHt9CLNZ+hGqVKMmR3K76Y5PlB8Fq
L6bImUWIG+oFEZhu0OPzWTDxtkmfl3ke5C6jhkOn+pZeKYLGSsSxi6UtMjopW4DIZjt54JqLVa5i
//b+6Qxe4GHoKDX7ECC1oYVNumYxeTG70gBX+ateEy+D4htf9PHHj7motUnfJLUgoox8Gu0xdt6f
69ZXXnZ0t14Hm05yOlb7A/9aYE+wQvE6hVRptfIW9RI2gNz1zQsxQCRr99XOC5n0u+iowEsvXVhC
+aS+Mx6EaRF1UFTAUi6Mt6fli6xbC0/Y3L5AphfEU8kx+h356gNAtIqaHS5nrEQegV9+gIAFHaos
ORSJaAVcCiTTEJT+h/NBbNSPfB6ql6Y4R8mW5L8WVJj9bSgi+JVwIRKdsvmBJk5z0cvSK0z/gkYE
b4zYcK4agXp6hxsh4FNjDV+wZxbnfl6xIxxHMAFpv5gMcPDzBS/INsQvjnIlJ2ry/fiuaHte/Wn7
N3pl5plWYpVALsxoOXWfeSfO+eukHOZkIxaZIjlXlQxFVEUs9gmEgge97r/eSXLSxrNklSS0SfzM
n38zXxTCDEHzPt7C2BJScvnOcyc/tvvB7HpRIBRfEfIjmAnOGA6MsfCi2vzqFuEvYFf5oKLAspqp
NhrF2NAGkEphyxXrc3bWOjvmR8FFwoyfuE2wXYriIPOsBpTZlXlSY7AuWZJNol6QSvcl15PJcwcj
LiAQNBnIsH6BvGTP4HG/ZLhE7hBYKgDR4tfdRMALxqVQinLIGoMSdfqKs8OYnEIiU0tYTNKvCUeu
ZOu7oDkzrVWJ/YUGTvr06jgLm/Bu2ho44Rvgm0HragclupR1x485noaem8C4FTKu3ucucXVuCnmL
M7gEaNjHUBbx14aPm91EU+CiuetJ2OphCXTT+L6bNmLv56cu++p6pIO+I6GVJFdMXrgJKHotSZU+
3PJme1zYedWraE/iO6npILKcmrGEiV/VRUh30YXBURzHW+3zs2de3b1+pBfwrEDh7gnZBfWUyil5
GsJvZdTc85YlOybdOAVnyUCjH/NzSRlFITZwCu/9tdNlE+Ye38cMLzGOCTLJAAaGozhMetLNfYUC
tEGgUqgmpcj39yvhgMNG1CqeMaf0sQ2/rKKDOtvSsiS2wu+aLhG8hvcQmxohb2LrZwQBfwOjB4tb
EII1xhoNJAlqlzGM72qe6xDLReRY/A9kqMA+6tRFiiPOFKDcyXeVDEckJ2JtvZJx1+8Q921KA+8H
o4aZXtDaPfwXGl1N2uReL0Ua8P4F2/AgjRRWTzBZYktU5xG8eaODR6oZxFBqPIudq0cBGtg9wn9z
MPZop8cJb3LAj0yA3VYiGF49YdjfOzsHG3MeM5cGx5968keIi8Ttz6mtjlU8QZYumwunKfngGemc
cnUYYDXr0EmkzT9M8xUzYn31RytAL/lx95FDGsIwfmrMGqDjsJdP4VzToUMVqSWEc2lDqIMN8hGo
yJjqyX0cRMeGW1mSsvoev31dV78SK0R8ptNL2D6p/7thGRN+L74TF9udwz9lDrjfYf/JmSEeZn5n
P7SvD8jtfyqS1thaW4BworcwB87Ez8e0chytEW3ZVFErwCC1JbkTpquBw3g8r8hwKRo+FzG4rF6Y
qa44jnQJgfFc+IIsqzeEU/m/kPpth0KZ5N6s5GGooRe2YUlDOYdGzqIti+qvpXhf0z+WL3kr39ot
0Ef9933jnzqw+SRoD+9052h1W1ZsbBICXajW2DfK5PDPvRTdKVB85tsYvcHEHSU71wLVM9+ip33I
rahjFP6myAhqu0LyyiXqNjG1aBjaHy5FFNSR8uKIjVgt8E5PWAJ5BdbEYw8PWK1lHn6vJvVdN0Y2
preB5r74O3NkrQ9jrOjFdehbxoO7SV6WXPGXqhqztQkG4I3up0aUWV3SrdwYwT1XVMM5a0L1hiGV
6oVfqVi86nleFDXCi6Hejs6/9H+Wnv1Ol/5folZfnjrvE0zvdop6YDWO+1XkgydpcBmmH3uCJyqM
gAh9a9P7xpfqvYliaYc88XA/ahS3P42tuk+KvycjcIFt2EN/N/xLseZX8MJXmuYKmGwFfDnJKzC6
xmmEHZmf32q704P5RnSe7zeMPGda+oilu2bQjd2dB/W0LV/ryk6bHEzgga8STCIoRh8lqwU+3Vus
EhScMWf3R/fEfFqbK4h0xnPbRGga6lNCEHu7VY95ZDU5VZV/BL/AgbupYLYy5gV0QF4PBWi+5WxC
zyKiiOoxIUDif5PWKriGMXRQ2JHmBO1vfB2MmbdFjQnXaGR3ENQ8LzKQuZhXlMY6VzQM1oCQ9dVj
Z90wDbRUqKn3ABXRsxARDdb8H28wN6MP++ciM8RszPDGqktPk9FLNT+OBoHiCBnzIBxM2PFCRBmQ
4RKPBN9pqFk3rNyJyviZuKbwKiz7aEMLvFAoKZasyLZG52Qkf6H12J8UKRyBPoyspkhPdoAi/3KM
vNWnzLR1VS1pRtZXSajLQ79J4XUOVaZ2T5fe9MAPo3txSnhZtUrQdCINRoVycEihoc7fBM13dO6i
qGP+WbeM2J9exe3N4HD5NMbDSiSHCzEGDbsS2CWA2tDlO0SQ8es2xNTBIGqkxjjbSJxOsIRzR1cS
NmGT+PpSc6WEgkHcJvgQTC9Ju65h9x6OpUy8ACBrZDpDCHfW9eJ5+NkCQAZLiFMuxSVul1XUtZZs
B+N3grCXEvSfjJqyEiY+L7wY3oxYHs3N7aFdj7mv86rbPOUxf2+gtdUUeOFac1ZIZuCtzQnjAaYA
0xfuhZDiIymBWd9siblrRhRUkkm19G7SwJGKaThFsADDi+y7Pt5nlFA6fbCvqIaGHnDc9gdmOh0p
QB2swZXuPnFNxO/Q5NuuzD+M2Ir5qbO6cts70trghgqeNczjG/CjTEqGbvBoz9yrHwjtI0lvYMsb
DTOfrOztqymj7LLSZCGN0ENu+kKZTT+ZX0jtZWlBm/aanC3suNjDKs+SiWdZkUwsFAgu3GTgO/HV
fEjfo+oNtsLPYdM0ZhHrpJ88f8EdwAAkARrKncWZtJVTg3JYy4UCVssrIJxFqWmfkBQkHbzHTEOJ
IbayDpVd731fFJx5u2cDbPVdDAEzad1VkdcUD6gYB+bIbgR4egHb73d4AakOOiR22SkcfB62r2U3
Kf4o3jXIhXWxqSF2zn8FriexX4GaIxFORKB+XyuGDVnXARjsqajKotrw7YzhOqcuMxVohZE00Oez
3e1N4b6ejOPrC8U6crd6BM0dj1xPtharE0ZZrmsH8kY9R0hh8P6iAIdv6K518D4d1eb+UdLa2BJF
0X23dSciZMugJbaAYqI7INzGu06dr9DP/eZRE1TCbWcbUvgIvs5Tx4QeTdyM8wwZOUmJhjFWAWaA
QrDJVWYvAlzlKC8zTFkklCce5N3Mzc7sBUiUHzWkqYFN3BIb8Zu3Of26n58KTzWSn9OPX9C2WPKq
1HEvX3MjAITilvQeqeTRKaiD4D5R/AwrwBrfzFPNMT6d21a77FGoIaj2lcZoOP7Omz7hlFbGgAx3
dqpZ4iVm1sd3t+onD2zZVW824NdK85eGVSErmRT2BMPR+X/1gncp5tm6Y6crwqoeOdkQCZhWSwNH
YKd7KSViPSXApoGhM1tpGt0uc1jBL1Ri20BEv9mzdcweq+383AnQwkfo0M5VFAb892g2pYVSBUAM
wY3NK9lJi9ZXOhUfVycfZFoUgJYN4SLKSmWnvrQuk8w/OtlmjhOv8PWXvi8L4FKXYXG2pxvlasuD
+G0A5a3dlQKDRPigrgFzoWCzSRdoFfV4JL18+HgIsgMKByO8itPJfd2e61c0ywbYPlFkeLbyV06M
8waPoKxS8aB1g8/QWybEDn7SzdP1nC6YiSemBj71Oli/s29B8+rqalIkmNQnK9bdt1BZ+UdYz/9K
47DROj7PXVbYpP6JCfd7UwrqoIYFl6ACAoe6JnIdviwiGTfokIyEZPzR3AmS0p+evj/RRkcNVIhm
EH+StpaljUuJ+HzA1MBh8VR7r1nlk6qVKpMflmUPqVeJRGN+598zZEQhoh1covh0H61MoOdknSmJ
jMgm4/GuEkJnX7scp4SVx1mdJk1bg3n3qAvJlJD/QFnR0Cr3qYxhxqQhnJL+iQ4LZ848WqjbnWs/
5fIVENhfUfBaveO1+f2GEvMx06dBr3zF7RDKpjkVMw6A2NlBeHzEhAYaM4hGCtrV//d4nProzF3k
v4kgnvTd2DNTxAkgiWMnZPauWjLZLz/hvGzwJPg63QLaclIBRplb4vBMUZTOdB5BLjDPufhbkMhU
haXxlni3PvfQoU/ba3Roq9ikqBJXId8y71e/Z1Hk2kJQ4GErrc5HFJueitaD/hv85A1X+VQCHlHR
N/ynhGs2ZgD9PnMwQhpVwMAnlE+3SWWJ4t0abihU5C5x7IF1EFlMqHf4jnQBTRGHRVJH7odZNP52
WDBCyHqLVCdQ7uGQ/MSr9fyV5EDps2UAfwk7CuIV8gMLe149xinD0Y9aCJJbrI4NMmk4QhHPBZoA
FzPDGvR4sYEkQe35i2mHLkmCd1kEXWTUKcB6v6bJClQCVHAtP0YeUiR0x3Dme6Ch5zUvoy6XePi+
k7Aq2vEQrael23Oxzpym51Ip3I4V5vDYmn+zKmRzyLVIXgTm//O0TzVPp8bXMZmcFss7VO4eKQc8
qoX2HgdiBatYCUrFmRdzBDDlxqNCU+l7FgcUn4LxUfCI8SaZw7ZsePZn+UmrAFBjCarOtDH3K1kp
W9YcTcRFc0sRIsdztvccIBX4GUc7PUn0Z6TqPuEXV1WotCPngLsfTom8Vx/ozzqfGcB5DdvYB8fi
6tJ3HF7K9TUqYjrU/OmmolJsqXKBj+3jYfkGccVsbPatpExbpWa3SMdZWq1hHYwFdaoHPg04OrP5
os+Vh3FSjFSkUZW3ZeRIj/HpsPbzVAAdmGzPLYt4MNaPO62jrqB+0EkgC+NOvp8iNSYBNGn9MxDm
tcKFwNkj8pnszfewe90nZMrLfLGHPP1dI/piFneboYYIlVYhBsgiwp2jycofMIkC/V6mxfMYP3fW
33NF6lv2H0da1qwMV6uCNpMviWymv2polnatPulUnUkDRp4igLTJFPRwfggThe4oF0UYYDRDgEJB
gGcRpC0gT9mK6ZR34jAqW6TMkdS7OLOfxAkDFBGjmeb8g1k5fr+G5AaMQ8Zz5Fawz5iciacrZ67s
WbFv6jXm/Py8lkxwQ3c77FW3efGJlgIIzzbR2azDOnI/BStpx1s6+ZQk2uzZ0dZSS8btAjzj5BNz
MSzbcI0/q3ILRX0prRw7o1MV+FmtjDpa3Wmh6vCqc8sT5tui4zVEVx6B4NR5xD5bmh7jIHftrccl
6qjUoZ9is5CwU3Nre46tkPoIMH+HpibxCzAdx/oFBXFoSMK9a9U1GY04CURYTw245/dQKvaaWh6g
Wdhm7daonyndWEl59pEE851NNJqXdunsLPfouLHffUfqkcNNFAE2WGnd1RYsVkhLKWmplrh5n+Tq
2KNs7UyE0l9aPSOBBM9CTD6tehpoxqT1dk+7MrqsIdFttJ6jjoQjQvsJSRcpkKrvee+/oyNXaBPw
4GXfgdJYZmVKn4EZ2Zv3jZazIAus534M/UGeP1sjvtCi3KIK7xVISfE2eBvCuZjPeFFIFC6RBjp8
twFs1SLxhWvkUTDTLrNnuwaRuZe3IllVJVJsV9HcIR13pzPYCplDdO+oep8+JWML/enN+kOw8tyv
pQt0fNTnuZF4eTzFsttJy9q1eexIOqqoDmFxHfMJW2FMR1bAZyd7AXWmZeqwav6FYd1I3HvUXKdg
+9Finn6eOApmKEuIci1yNCgukQ4wx75OceOwSb0OchoLCSW/E6EZwgfzAc57LWhN2fiLXYl9/gpd
od4i58JBRfpCfDnOPIUGS4YYKHgOdpfsx0FXg33CF+lGeRZlGSDKLg3XQnL34ExdEY3SbblSN9hI
4ZdXIWHTsQ6nM1YR0QLNLkrAguhANPBfxpuVzS3ozaAP//eI3n295zLyrOktGRXh2mcFAjlCfbSh
mc2qFbIvve8S5WgVQM3/3jt850WRUwYAve9jcZqSSdIPhcIaM5nLl0NK84DuFkXZS94cmaolY5JF
/tLEuwL6yxDdVDy2sCe4UwtD9LJ/GeJWYMUJ3PUId3HAB3SLYBqTXFNWsDH8AB3hrrS2f7rBqxlM
mGEn0OYYWxVW0KWqVMTMKsjbQGd87Z6+y62JIYVeBwdP+pO3g6kt/pkyRuZ/Df2u12yDK7yUT66z
QaBOtPRY5kZB/B84cKpd8pdFc7i7TY9Qb/pXU7uv03ymsiMHrVYNAp4oNY5BzusQ192octfX5fJX
2BKshjkkF8PEbq7GLeZLx+spIM6rP6cMqeBOH9LID5I8lw59DdOdUlu/eC0/tVZDx8wILBlxrBvp
vhaso5Bv2qjJ8Ktdq/J5TfnAmBwYMmo2YHBSoDK3p3qESaxU97DrOQxWtQmpM+7mx1qMqhVTI16Z
fo50lz0E6DOjjQeqj7eDcDPQ0sdganiNqE0bSzxgGIxtBGs9hLN0NrEBxBUqf0gyabWggOqUzf25
19SZUlOKuJ6BIw8foD0HKDfEsWLHpccp4+GCDpaZi+c7NPTOO7vHd3BIimi3KeaEjkxcZCJfMQJc
hXv2xVXpzValG8+7TPQ6zpm9A9YbtPuLSeDMIas0E+vSFvMpU7XFmaeDj+gwwM4UTxQww1mS8QNF
P1l+MYmjRvKMwPGCi6Qxkhzlz0iBR0uFsvPtMtBAVddOHfbwVJokB589iUK3JzC1cK+s4vt6uxOW
2rdA4h6bxjD3S7htDL6uyFMlWI3E3WpBp5xugPZK7OyvnTbygci/EDHAD9cKaUrGsjLaqWM0YJ0T
JPmoLYcV7IG3cSTwFgv6FdaPqVVTQbDzHofig1mEfE27IpSEgDfJzoDl1kh9Yt9a3wchvKEs8cwe
2bi3mqrGzw0wVnCSkXfn1T1pnHqzayRX7Tt3D/2t0g01tyDXF797axltE9ssQiUGzaIYsmdyFsNl
0loQ44zZWMkpcjazEFXaSfYNDZMYPZBHibV0rL6O0P/TqAuegB08xRL3XWFPUcgDjve14+pSTEUR
jTA2D6bVkklkWvkEHCRR7DAM+nmXcMfQXZyBF9dEQVGUYwaJSNNVpHdZVpQbOviLBdY3pGCBvcRr
9LWSbzhG4lXTR80NrSvoq/XfiulUvnSUS9V3AxbE927prmdLeGSUK0NEQMUQHF+uh5sLYiWBwJbV
sPTglFUv0xFDcQfxR18ZbiWtbD5nU5WX/P4kVVvPKP+oRw/E0sjXYNLgOMmHXJB6y3s1/yMkBtLY
EI5QKr3bg7di9OqKr2oFYrHFw+4nFTrKw4aUXVOJV1ZeRicJKlc4/sE2alY5UeQDIlkGrBzRlqHt
YoeWkOqrgFStcF36Tkekxk1W+oCmwdPbaPJO3zYWesGBMmvh5CWldorjQOh8NC/ViTSOcZaiNAQA
ekdLHFMQZ0KqVMLAESgazJlTrwlKczt1bS1GAHQDKCC04N1PQDg/7TNbsy8p+HK3CtDifBxJqjtL
ocnpZ+sl6mkCtHlVikLrDEPI5XgdN2oU6Jt9AupIUaLBFz5vyC+t4CfXgXq8u8js6CksNjRu8aeY
DcW+QM8Khq8azJP/RQAZybBD/NRxe43ret2afBqcDdKIWi336cWLf8xS7AlTTe8G6RbGdPUOL9JA
PejOB4GqjKFUGRGHjYoSuXnnnrBrTUPjP1UZFpGUDuD3Xx0oBuqU+WPCls9jK3bBwxpqld2oNZNc
nzvhoz6j7Q0XKWiQiOHMHSm9YoIXcOrh0BED4Hy30zX07eUnEbVzOh7S1ZRrUKTnRXfIlvB/4SaA
oAkeNbtqdkeGt5XFkeYK0HN+ZjDLnaxB3HicLKR6UMxPsIpEShg7Jx0Ix/hhojdp7xbkBLG/X8V9
7Or1BVxe3/buRBhs6UZlCwk1A6v54P5LFOzMls/0EeWIfkVU15BhLTdr5krCiWMmJTKSSHZpCnil
wL508AH5fmK9xibiLkhm8gCLSYLMDZD10RPCSkPVXYpiS8uBWER5sa8lzZ8EDfEdBTHRqSBplx6o
WgL77ZTI1C/h//H7SgDIPWSD++iaJLVt/ac2jNcdogh61/rB23EtNu/hUo5vwxJs9sQk2MjwwxYl
UaHNGZS0HGAKlRpgUpNIrQH8DzE1pPA/pHz3RyjsQ+2BJZ7RontSPNqE9doUPuswc997x6tWhfN6
/0k8BI5B9zpr94eq+ouCNYmIzJVzEFnBhbU2Fvy5zv3aJzj7B/qF/IMFCjMU6g2Gmu7RzdY3v2UD
rISx4sUZbi8JpbkInU/sAmqVjQAHC/GJg92834JIqCIYq9fZ6qK6iDLJva3tiRADDb+BHnPh5grL
TeNIqvKuuFE54xKHwX5dVF7m1gBTRKpiE2WQLoxkskZm2+jg+ct3fgwPPYjQg44bDVofpoXDZokS
1kMI+umw4wfzlL37RmXYDeIC83Ji7qj1x61RzmPNpIKO3MwCos6lqjvRWO67ScreyshqYabvJ7sF
ar2/3ndMSyIJoFzy0CzbMRqszG/jI3V8EGjZ+b3AJ5i3NHdmxwFzH0KKVxysejPY3GAl65wWa7yk
Kzu1RtSE/W+OimFraAnqGhuuB3WRbmn+sFMJtcoGh9LTdwMRLKqhl0XYpFwxa2bi20L8NPocpmxS
rNF4aeJuovj75PnVwfg7ukL1AMFKxlnjDKjq+9Zd/k3g1sdKH7yPxjweK57krNuQIO/PsUvaMKql
STAJg4P7C24Ip/fj87tyscb5mDMr1CNDQZJpJsIY5MVNI9Ww/oBUvYRPVglUXnY9Gl7G3VO6feK0
OOq0yZw6kcHh8n7MJem045XLvP0UuElYXCicR0MbENVFb87z9wDT5gmZJj3m14ytnW8nG14jRK4X
6ukNTZcZNw9xsbKXkaiVOin3ZHMPVnfBDdZL7MaCmn/fo7uh7VY0wdQ6XZLj80bxZA5tL+/Dx+Td
twQnGkMa70gubFULcNUZyUrU4PYOiYk532SVJ02RxIJxA6oCy6ebOIwi0PaXXraxNnR+LftC6tbH
ondG0DkBJSMCSOJwrtrfDTrjv01+Lnzv6f4XwNU0BNwrEj197fkmqWmLrPcJQPaZXCVmdAa2wS8e
hmkr14hi/zFhlShJtafoJVxtNvvB+sfx09pB0AuWKNZqzDHb3M9OnMiR7huUp8EzKU/FYkt/HoSZ
G7Cd//uR/+ls8FkHZlvEnT+mwnG8S1DSkgw2QOmNlXwS5zQilYbM+z/Cqa5DrtDHJ0ws0V94/m1J
NdtdSawIbkBbaKaFS0SKn0XjE2CjYAP3pd4r5xEIXkMya8JEbT6TYEuB7rgkdTZyWO4zVD1TPKih
EOS3yhFovIRHAAIBirpAfkpm58JrgCZ/Ns6vv7LJx4ULm3IxEkJsTytqkWDUCBGpj4sbq8DAHL4O
T1ArV/TbNnSKxxkPOIxAq4Wxg0VvuxNk98rxOawFNfIhfoeWOLUNlys+KxTUsOUdBj115p7f6HTv
jK1kQM2YMDe4W3NfIg+ow9XagRn5VosZ2OgPhQZu5kUnTZhb7GybFFFdX6S2uqOWVzuosQ4fpxXr
X8Pp2QeGa5xYUZO+2+u5oOPakIiCRloijw4TaCRSMkbU9s9PJfdR/LAQOlC8DSoXv/nNrXnMY6VH
mvYjIf7j45j5UnRR8u6Se9nQ7B6ediiO0CON64FmN5qS9his8UIeZcqecG/3giES2CmdCuEor0lp
xelq0gu9MteTax1NPYQxzURzLn5gB1PNCmybISLpbnVNb78qEuo1J07FHCSuOwp9o/nJvufqpV5c
xYVJ1wb+T1r0Kh4I7ZK4bUxPyoM/ntoLlHheq5vKEX4e1OV3R4VrucUt+aYnHPuS1IGI+RI3pZWT
iYCucjLah4LE5v3m5CHFX6epfWoYV9dXSToXixOXlfi84m21XsB1lYKJbG8te0mrJd/6qlOWxzo1
yx81LGaiTE3MEgPeaOSPOevGYyGHzaJ+faVRgxumESw0IwX68t4hOSmSCUeXHKPPRy5uUBy7Ga1P
99/JUjpEL7MnBQquYeHVcHcQtsELJHRoHEpivnhPMnmB3bBixB5WZKgNc0uh2tgF0QuYmppxboMH
Q/dLkV1HfQPymTU5g6ZrGKK1XGCpYdAdz6efKv5jf6aQMERauGz9/W/YthsX+M+hNd0fRteOM8rb
N53HS5lpbVfmyIG8ajZZbUBOZlXnwS1CaJuZ9F3cJrtPWjZPfGONR+wVb7hBcLHi/j8L0HK70GGY
mhGXnvSZCKX3f07dNRyvk/JhXPYgCLjvVlUXCo1SPxL9+GskErmVb2h+LVv9a90/E/vqXQs2Rf3G
wui8tPltpBVaF2ExUruerq+x7tez1JHK0a8uXBOkvhpQYNix9sRiaHQXJvISPByoWC5/KRjzUuPD
fV/3ySGz1JSrZC2F0VT7eMk8gkDbxv68BtthuNTLMwa/dUfv09R2HgRIOYY4lyWaN11NGYSF/apk
u0tJcrwTOrXqEuSVcMxYDSZUuMYlkczrZkxwwubfYSP39lGQeCTAY/DBkyJ+2TMxw/Id+5wQS8Xz
squkchKYYtZjdj6SRc3zKnvi0Fdd8ln/8TPsZLlkrXLtZnXJPizkelt2oIgWKXsDyw3SXFA1Dvgj
fyWedDKhK9bFQBtZqlcx56AV+Jani50Wq79F2LG8q6XX4qu7G53AyrtjsWFWYZ+wKw2k/m9O/DtK
DvJJVN1u4tIKuesU+Q5kACgUvVovAYRXbdXkdt0AF2A22brL1mr6+/d/YVdtOxnNa86uF8MIfehM
GFf6biwmMKNB+y9yh9WtzMt0r95xV6zzB2QV7XbmbudBezKSDcw7XKZmeBoT+mDOnn/Hu8u0aViF
LJHXitnLcIwSJI3BOYbRJSNTTQ/Z7Lzn5+m1UdMoC3VzunJuNvKEZu4bfJ8t22HYh24LVocc4qNZ
ZPC7p2riffI67dbTEelJEf6ywhqThlsj1nD5GIEAEH1z7ETeCuZVqeWnz5hcSqgSIyHAqsIWVGtS
Vy43mQ8JrjF9NR/sO5VdZQKBJJ/uXbEyW4pJzN/Ed+ITKI/16Y4GoOj4rY4VFCaXCtv9WWPUrr6y
+MLh9mPM97YivoDhU+cwR+c242dKaqKPr060Le48LZpr0XMiELi1/7994igELtezCcFZsqvps1gM
rektI49W/UHhb7kgpJ9veJmcR51dv7rNk6jBEwQ4GEjNKTJYaZE2WfOlTCIaGh2MiUsVspoWygyi
hIoZtQXiwgA1VWaSOCU5Dbf7m0EhnlEedy42vlGA5H8zsNOmTT40CSNnefT/q4dBYbJ0wzuRpR0i
o4OornRlqBTqZ2eZ11hBj09bygBP1VS/GNeXDwlZYf+TkkFaa/TzUuUdDhbje+Xn2dNCkwXJyigH
nHQyCbVKSxleJJ3xE32tDnNSDifKkek4QTRuhfEoQY20poUybZWlZkg+ScrEC5sEms80rID21Wq5
V9kKUAm6b/g7cKNggsz4mw02zBRjdHgGjuWkh7ZX8CGZGNNgwx3SKMxZ3XQe2pXOBNCf7j8/zH++
9ZBO2o6kheeTZsEATIS+xkQNr4hRClFiSIFjFqxn+VoLsFSi8mF+rn3Sq5j9Uzhz8d5kz2/lxibT
ESETiQBbQ8jn1z7D9GA+MtIg5cH8XNwumAzED7YwLa9aQtvG2qx+69U1W5jy2QdUXIwWNNb8bPBv
A1FlOfogmLKFdmD7KXruIQP+7yRdSMaiD2eDq+s5fRpbQoPhvwS9QeC+6A1LJRUh8tpJpls4SIjJ
Tx/KAicvLtBn5Acb1Wa+rTorLt7D/dmgI700xF5ze++h03VAflYxceVHs5PGjG3hi8wv/C7+rG+n
WZ+z9pYov9qj5VOW2HYbQSPz8vPq/wM2JsG9owmxWeqHrYJ896xJV1Xs57LFm8xR7LvTp8YSl1op
EkV7RrUJP/1FbVa4aZTdpx6MI0Y9KZEpRrtrTH8E270ijyyUJMIehZv/oTw6CfNBlPGMqJWuMgaV
L5bDNk1cNh6Y/XEMpho1JDTJRMVdWHryWuB2m6dz+pN+WbfPZpcj3wnHN7rRdIan2dt9xJ38Dtg5
7bqKEg5BdP6OOLzlCf7rZRryhjO5WOaMzT3M7tXWkQE6Y8F2I7vbhPp47Fm+2HeHnvzw89UPwO85
qeP6lsIJuRij6BzJiOhk3xb+KijpJ6GH1p0Rc066oKoLkZtCY0nf5KPajTfnJvoC0MQsdpCAC9rE
tPNH0YXgKaBqTma5kTRVWi5RbihmoZcVro/CcwEymX3kOhyQ07byDCfnII4gOsEW+sDRKJJ7lYr8
9T89GBAvOWF/RMYmblMd4ut5XBPA9aturExrH9hRup6DehvFcwgcwtpfJuIIZIO08BjXwIu2Cc9T
WR2PdvSdfwHg0NUaGHIxjAOkIrttiMommiATvRpWIKWaTkcmkNA7SUV4VRUiSSEnXOrHsnlJs+28
zBl4rNJ3FP6kgWGaTY3GH4YKUDBQpOSra4juRGx8fxIYlWluM3toSuvR4ATcZXMrpsf8PM2JOFOk
U9l5lZzkaCVYQZpt3MkurzVTJ1ToI5Omz7gjE4TZ8tuwemp5FMqdqeVLatyh0rUAtZxFUbF2c/UY
JLK4bzgPiy7p/Jl+2h9r3k0UqG6tEgl4VJSsBwfR2yrln1gcEfnnd+rhDtcEiVgoDPFy0AaifAP7
/cp2KtkNnB8+XpPt+E8pJ07BJAntg959V+RvzhDCTDpvJjP/cNu5iRKGM+tC1P0V55BdZJPC4uAI
WRJAaR0BcxPyyUfn/zgvP7d0MOsEJ9PXF7JhEkE7Va0AyCRkdzgxvS6IGGQbDoNwcYTHJ+HXZ55/
18bGOYYgNstWnB81PrhmwDeP/2kzDuMqviL9FMrUrsAmAOk2TipnVuiBsqRkzjsXCPLKNrMK+x61
tWs8iaZ+6qqKoefqHe/JjJWOIosItZLfh0xTIwK2TbSdQAhyDCUExCzp84wDCC3DSoEdwcZ1XAOC
JnSl9pVoZhHX2+O2mtIBKN+d+nLBXjbxm+MJAfwLWtwHuCJoK9hB94viQQrQKLac5bKGwTvErp0L
HznAQODOKH/6RoqdJpdFEGt5O+txgdfIPkIXaNpeeVRkm3E9ZtqLi7Csx6ohnFabp5r4ldqYTt7C
vP12vKJ61MCHPUhBfskCskTvmpoU0qCSRtctWCaOjCec+/30ov8hVH2XuZ+HtksQQXACbZfN9Kd+
xeuzCKRd9SjTRB9venjgPZP6aOu95glHreOv7ycPvbIPAxdrgxEKukO3w831CtnpkN0kHqLvzHUP
hNjOqOtj4FbzX750TZdrn24pWphcZt3LnCKdz0/kDlD6de0YgusYDonAFDkgjEMSMMLS+LF2Is8K
K8uBHSRbgSPzrP/isZw7uO+UXwFGYxvqOaSk2lyXGanEss+MXq6uM2WU81xE1R/WWqa/zFjKTlNs
cCFmfEVnrTFWUoEBWvoAFm6LU4mVhXL8KOw29Ar14sE6rQkYcM3HM4mQ3Ij65gK9oX6rhYr0aiqK
C7EV+jlM6pXBYA9V0XG2EEUYXXHninwb9rCh40g8b5nI1lyj2N01C1s1M9bzFwA3bUBu6ymv9LPN
sEH5WPdRMOeG+n71WJily8MO5GChnyJgLxGdZtKj052BkBmSYr4IdqbgPHyN0P9LIEfLVhiOd0dE
cyCOIFEwW93ACZJQDmQZ+Rud+FcRJYVai5F3eM1/zP5UdSvh3SdUbDSnPg+kL2K+O4cAL91HUBhO
iVXyiGinSro5cpxQuYP0XAFSV/Cs5oNI/YT/bkxyJg58CDXm54UZikpcwCiS5LALlBljcLnD8tDR
pY1H3rqSMbMwyo3Ty0eB3y4qQySQ7LRT3USfrA1B12aF0Mb7jrF+x3A8ThwAwWe8VhWipCA3gQdR
B3AhD/m27bahEO57RptNre8KxEMROa6NQhLzIVSzsJYQ0HdhJ8Zx3T9u0YXJ6fAnVO39dg01A4+C
Lhv0AO4lm1eUOLm3Vqo3l3CbTpgS1+uDHPrI7a71OIk+J3ZZGsOFZCFPMwbzJ0BCphR7YYgCIuB/
ELD4dzslPRYbVdClMEVAwQfDx5tXZkdx1RTIO2rUGZYn8otwxOmG8ZWlJ890vJc71rlclMOlIRn4
yEMS1GJMgroT17DbbrDvm3LdwqV1UkW3drhKAHDLDUSoXQPwLUcZvlZH5hd+Ce43WJo/L4ugRJAU
6tGATA7PYj1PokhD2EekHmnyuOMRDP/kMmNrB1fzrZJJAZQj5uWBOeTcuCgBaFx2AyLtj+8Wcsvc
wU9rg6Q9HQ8dskYtphx1WdexnLFQJexLdc9J3vZCZ94W14OTR39nin9h8k5tBOxxvl3O/uPvtKKN
4QtgFVXsf7OKJt50JzePx2zMZgb8YFmI65pFmGVh/CNRyJTis/Rp1w3q3RqF4eRATJ2EbJVXspjt
S46iaOXtDdj0EgGUi5MNKNmDwEyIdRXgBnYYVzy4F2Ht0rHALoxc1yMmkiImUZUjQsPNzMXIIGSr
ZU6qCS5E9P/wFFQzy88sBzIpWq0ybjW7555Ueb7HHMWzwqm+wCTZKQNNswgL9wfasodqOkKCbYSC
LUe91IHjNtP5YFYECt89wTVvFZcorSoTfooPP7+ZRg8v0nBrJ4poxfcURLp9guerQqPdYv9+jbzL
A6YnOfDeYZ7QvfIj6s52i/titGaFjEtaY1rgSw1Eulevfb3sUaDdbljSkc0nOQtZ3Q1paEAxOYai
5rebSzAdselJwMOTOwsbrDbrk2TF1RtuiW6rMBJWnwmr4i/WGvrqoWsexpnteE1EXciFm1QgpYJD
DAXuyrtIPmo3AF8a/W55DipOm2mZSxsm7mioAM1QuO7CVUsMwzqnS+XyeM6E+mceaXQUgk+birMR
wPirEpFyqF2p4t/4jJojiSwXGxMzopCgnd7UlB/0OWdUWi5LdijJ6rCDxhVQNrHkjuSBiHQqfeFR
q2eYBR3BfXUQQdSv4w4SPQykUhJ4fkw0jtL9oHvDmliYb6LCTMB/FrounZlgtt4comKqTvLY4dhr
/OnaNWLrNXJXf90/Auwr02CmlIGMhwHcs2NhkmJsPPFqDoSjfurfoEAu5MPuBdEdEBLv/EL3EMlT
SNtyfUaMl6G17ZghPOCLv1WfWN5ZNaAfocW/PQEgGbG4nEpMqt2JVTzbnRwuhRmrZmqDw9Ew5enm
xQLTeTje5qzhBq1Rm/5mFgcOc9iGt+o37s8h9qv0i++1YRbCw6N4QeZXnURcWql7ME+2pYbgBfhp
Vljn76GFrEtTXnbCncKB1TrxVP2Afj0pSmSvTO2O7j45KITH0JYL/FIVD0ovkgh27CtBAAKd8AIf
r6hjNWN4PnnrgSG2JrX9NXXjoSlCiAMP4GzgRfWofG0AUKs4/z+hyaDONahm9Q5MEEcvEosUjT44
5bvy2FTQokSUIIMmoBJPbNWZcNen25BPdHZuVmkvfgVew8nLy+a8fudah6JXj+XyjyTFzwgHnSUx
JvqQ/qZF0tU/MvS+Ah8Wx6F3ZES634u8mJYGt70TDVqwb6QBRHnJA8W3AnUdyYlt/bw8Q8gptBM3
4mxcwkisjEK/yZzRE3HVo2G7bLfYkH1j8M3D9TccgiREDjZ4d2rA/6v11+g5GZd519q3iMAbuLtZ
FZNskbJjsM6+7+rU6/LmqHF6u1HRxK8iHJsW/Q1lRwD80y9RoP2I50bOc7ixsElAG+EoI2aizTAT
hY52V9eKJKOLQQswMCHZb4r+/OZg9UcZ6WWIeDClA0A5UrDxv81Ja3ReR6V3sqhsBIOP/393FH2g
G7UkbfFv1FVol98ge27zzgcN7ElgfEi43WT7iFN7m1J4ld4w3QEOkLkU7AI3RIZ5kL2AtloSNtf1
W1Bl94n/p2V2ew93uJASqYuwKvw17TycYCwjR6sZmcqEIZjJkQ2SNhSo6/4GBCEFEWrSG01ceKlw
FyK5G5YQB357GIdtcVcVO/lDttjStvK+kGyijt7FSc9BzP0p7cfDnCgIxJxs98R1MpIHZLBTBlGX
OhT/VsfkXBedwkUAFRxpAQaLuWJ4fs8+no3dGr4CSoS05lg7gl6+PLBctqe2PVYbTWj4HWOmL8E3
QefHKcyLN8tPG6RxxTUR+bJSgZbPjDFrEheFm8bsnubho3EeR18wiVRiIOXcsZ09xXwky6pzfSC2
NFc7E4OhiXjIJb/vh8f7ydcEPpJb2KgLBVC4Idz5xth9TFXNeEGKZ3UjAg6W2ipbFg8kfVuNvZX8
H6Vrkiw0Aa7qhs2O1DmaL2V8lUurT6eYdXoGWW0LRZmYipX9QvmJykVydRH8Qw2rLdhXBRfpNnW7
P8eMJ9CrcoEs7UaibwyE1A0j9QrQaWL5L0iUqFElYxiopzuUCeN59XJWe9k+I/jG1WHZVMoSVy4f
Ldf3Rq7/xDKaCKbIyPEXQ7yKGzdI+P5UR6aEJMCKCld+mTsws/Wt73K537otG6qzj9fCw6W/iqED
kaEASnAO6Mt6qSBrgginztnllqOMZbyE6RI/t/iFUM4uPt4SRC0Ye0aM2Qq6ypcu8H3xPEYEfYJA
+iKNFdC7cMGSqaXJ92aRn370RCUlcN6CwJEljVCULbYNfXkt/DovkDFV8BPouKYp2EybV3Pfjp6C
fFq4lf50heJUrdMFfSEqEM/fzQNLnhwIWoIc5pRdz9m5f1a7FlO0emO50gMveYTz2qNt/nNe3STf
1xFY9ujityq07/eHM7DwznUcSV8VUdoMUSk/mOiAaMrVngIfeXPjdxNaMNVNruCJ76ta3fxdOudy
bR/KZfrStUrLeK2tY8al/Tn6NMhVKZahI3QVRwJo7lhfWZl74vXYQPIJBlqDDR1z4sZyrCt6Suh7
KldQz9GFLdT1TkoqVwE7oJ1YFZrLXLmwB1/StWITSnHc5qUyz2tZR9dA3joe4LYw+pg8DjJNTIdM
0MdwsRXOOVYiWIbKMl0l7uRrw7lIqLPJIEu8zR1yq6JOSdH9ug4IwUPdUBx52MlzplHaFsCZlpbe
9G6vbr9tKKo09uSh+7JW4zL7WWOms36eUgfCnkHIzUYKm7VubUPLGGMrw7lIGHyc2KafkJOB9stq
r2hZKOn1Fo2UGuJ9Nw1bYK5zRcixdCEoGB9VMi/3HVpyiWZXBzLiHo/uQ6Bi8dLyEgTzr+WhuAZp
qQLjXdpKzqNlCmesujxXR1yHfFpBppg80U1wFnDTS6hi/64sRBkVKcXXOiPcx9tdngXaE+ioRHY3
xrOeUTcoh1YhbI6kjWwjPIwbWr2aIh3h4rdiO5LqGRjsF5ks4nkGbRler1ZtyKiBfevBWnW1RKl0
zfOtpTEm4a/eBa0n5snvT/EhnahzTgN7uY6jn1yyBN3MkYzhst4pw4o6VP6ihGeg25qLsw9fRp6Y
PXVN8ajjtfV1plA6DDVyFdg4MrxRX5j50i03YTkK1CwBirgBHDJtqehgPturXw9grmPSLKGaZelo
iQuKjiZP6BcwNFvV4q5/VXmchsaizhCo65dHapmeQp+MJUbMo/qEgWg3mcWUDgVZoagAu21voUww
//XJZnArurwtSwXUqgqPT0qaYSN3al5vlQ4y/GAQbdKpDRz6l8aMpVd4UBgtjpw6+zYMe9COPN3p
kPLcKfgywWE6aWjCVfWXcoOEIVRcn/FXSUqyfLFthWg65gws5cTVtLFqgXXynDfQuBNnJ/jH9sSL
Fimvp71ccteKMB07xfgmJ85DbMqo8lVAd/7TFa19jCC6CwlzGFjI0uEdhLBkfpKHT94/aQLeX4BO
fBgqX4Ex5i5WHCLmbgg3+gbZvSWxZEp7kHhK3G6EUtebEPbktjUgE9i4nqkYKFlF8QDEkgEjeFEC
eOhQJtlODxUUSjR+b2MFkro0bnm4/eqmHUMkp8qmzGaY3rQ94eJNfaIHyglucr/Q1cRsmdmLUKPR
cihnV6ALOvP3QDqBIwYccaEHOmLH0wPmmBt5OSbOm57HrQUzjhI1gI9yItCejX4tOAy5P584Nc1J
ctuU8043LL+0/iHauEQ+5X/+MPXRo8b96BtPSYrdGDBqeIh6VJk5VDoQFCPbz12mTArywkuWg+IS
2ftl1cXS8FG1I2a2HVDMsXgpGuSeo9DktLh6pDYJTW350hgIf9cxb77EyfCsw7L6hi0Q9L37LD2y
BHjHCMGL3w5n62hRYf5e18T3j6CME3vOiJKqOodM4E1b3FCr7yo8PWmn460F7bJ0pOvgRK+BSma7
ZIdKSuJk3EmWLa8rObmVWzfKmbrOJinP1dlVMLxsJXIhFV2sYRz4yf/2MOw/8ZrhtRiDtEzMWBvQ
yoVikOFAaDyDKCF2WhQvLqZ/mA70lQ7ig+EJr00fsZMMgQHz5wR/WxjJoE/kZRyCOHvWwWQNWPT2
uitjl5zz3Yp1ao22tqOSMsFprys8a3yf3go41BC9WZJj9X8EhCWi++ipgUAmVcoqqTrpwrhwUvqO
3nNC18H3l6SbCuM4ahm8hkqC1ZMlvIoyUvvdIxkL6iK4mjAxaFQtqrhIfz4cep7s5eZ9uorbSGb/
Qt0CMhFZhXwd+CCfRuohxnpGStFEkZuYk3WfdSo/aOyIAXPx26O4rrMjKw+0h9T8oSo2XWnjUxHB
/9Sy7LccysV7kNygKI/sNPii+cQj5QYNebX5X0q847d44cE6J4nT19Felo9swmPcUlhUW/TOhHgC
Y6v0PtW0oxgirO1/lxSWE264v2zIpVTAvph+SMa4UuBzXvKGRNXf27SutMMaOkC1MLF82JqpRAwy
UCzRZKp6aF8Kcn+J5PvAckzVUAdKs4Whc2bofXPKNcvgOZDCTjtFTpC8OUK6zQZtwh+YhjJqw6Nu
CaweBBJHm1nTj0U24piGftZmpHoHYcxWmqemMgir++RWTwRNo4icraszxPxQhGABwYmaXAla/egm
kMuzcTdv+flgGcg1U9Hq5vHEWKvqCS1jrmF8NV6vVSOpI9Lb/I9Z6O/r0O6E5dbDM9oR81PiWDTa
Ag7qpSL72z4NSXkFCDquoH+K2WWyROBngLLpb2hPUnW823QLsMd+7WVWEYYYY+sjONi8JMmqyDN4
9zeYC4FwC0oHoyOK04SvfkN2g8Y1h9AySKKNG9sF6tNjm/MbbGXnr14Oo+tgy3aspompKay1P3lz
s0EC3IU84Nes49hzHwuhgpl0iNkc9THJ86hj6hPsXpRZ1ZIKaWTXqrLWxDBTd61vgWZNhSmLR54i
2hSwXRoMkXQPy8//pDCx+QHsPUpVUJZCXRhWcWe1kc/t/M0+7b1yb7hkgXWqs1MOTnJV52NY4Ry6
2SDTrRpVf75TlxjfBwueisPLtDsVhRu+O+1c+Y2te58fhT2+1UhoNY1dz59qP7h6OGUzwuWD/nyk
V5bp6HodP7i5Qc9wUT3qrFGgrcBz3kb+80NbZhcT5cWB2i4GvU2Y9YgoGosxOH5cyOloGkZdVT/K
Bd4W1TKNdg7fizHlyoV3tw9L/7K9N/hCZV4Tt8+o+chgp4n57YUHGcw29rtT3geIWiwNfDJWoRD5
mMZdMowHBrkLJgcSu9WUZe6uyQF5JmrZq+QqIebCk3ftf2G81QdZKbP3jF2YByADKVwwb/ecvRMo
M0JHiK6lNgOa3cuYX2DcTcAkRTJHd8HDwwWWcxxl+cUUgVzdp8m0yBCpbi2BhF/YZ2CmLPWZW59N
H/qI9xfZ0ZXp8ng5fBWLR3in8/eAfTcUYmv396AWyAbxntK7gTZF2R4KgiRvcYTY+jJKbaGoUA4U
KGMNWncPoeOfN3KgBwJx3veoh3uJsU6zz7x2OXxlH74P2Kg5QWN4y8ivlwORayUGQQ5Y+kVkjQIk
9QukesF4LvPcPEpS9RlW7MDMVegbI7QB+agN+ZNKs4lTP98lOmCuh104/fXGRlVLAB/8VM75gfBJ
49M6yw4gGfhvYiyRfU1/bQOz+b3WdxuTIQEbDTKCLxOtL2fUniMCQDzmt/qBCDaw/hvx9KC5JXO2
L+4VW7J9Q1gTLYmzqxMYSRmzLRzebYVRd4ZlnRUnh+nFFvhcZ3kUwrAjaNqP5mr6Rhzmtwc4aJZV
7itEm7jvOCP6dAhPbpfgp1r1jPIzRlUx0duasR1C07jkw2/iPUiEO/nYYlrMX0kK3M4noDvjHowi
iazRMPMfpwE7JP9QaQu83k4V4q0+eE/JntFKvNmRwMAZ7F4DDoSjsUGepHR2Zchv4F7Txk96KPuO
Hd4vve8HdMPIONsN/ADTaqV9/p0GK5iXcxnqZ+Vl5JHvfAiXJY1eHwvHe7lj1VYpuxQ1Gk62h343
Mx63oFkJf45sbWqU7rTzII5tNWI/nxAdLuxUZXyh1/FfPCE1XMg/mZS85fiWYBk9LIWuxhobWsq9
iwN7UekokKQljUwzygX8K62K5YX+EoErK1Ng+7tElq0wRMk44ljgUR3pKCpLF/nbMbZsVbsF+V6/
nkUsirClJMWf/vJtRq6OQ+AqKz2ZdVGlWtosJ+5E1MbBmcKIdz206qoB5k3zurwQtfMmhOPgikq7
IsoKXG+lSNjLhqSejphEWUAIuQsLEOKOMq8tNLdW9Wd8rgJNmQkdFwQOlBw2omasW3BNNCS3iiGI
6k+b3Qz5JbHocGRzfmCTLeoLXt1UtBBGUNB10+6Mc0ZAAHYABA/IqI75wConof/8jOIynW1A/A/7
vSlk+fr/JEmdDAI3r/6fhQjWLB2S+N0eAzjsVwt8dWdCp6RHGkrqBpzlkjYTIOxSQ/uZHfENIiNH
UGn+LZhSM+gth2KupnOXlHjRo7NnSZ2mZOIDGx6veOdOZ4GcvU5OPr2K70hrZObjvxdib60vrSoM
zCXwV0Lxr0KQYNIpSAv+1ZDY+MM7OMVTo9NZ8tEnvu4nzilksY31uZCGcVs2YmYE828ma/TxSiZf
iIKX/osCeCo/gSu7kZrfpaw9g0ORtsAWyGO5TyzlcJobk3nbnYbXUi3e8i1GGjcUI+1reYAyCqkx
YSC0IiXPoVVNzC+ViKEdOmk3I84MLL3jH5a68Q/9j8At/DXXgXbKMK6B+YxgiyMFc0s74qryM+Lo
lvF/96gh5PW3f0mOYFysQovP1Wr1tgckNXrE6EfNqXcBsy4AZfn6kVch6rqQy37JZJjR3uuUPcxR
4IkRAteu42l3MTDHf3hBL3H+umWrRkO2XqdxDEso7KnMELaeT7O4bDeTEoBfbsPevn9UAa3S90ia
NweRpsXtSzhALQdatjEGoxjTo5xsQmxD4GTklb7pMUI3SDGCcAUO+rZSy+hUt2CX55wgYKBVnav5
iw1oqNNOwmtFPQ8BuepJ3Yany/EyEQb0AQfnhmrQjQYeg9lV90FwLahkh35eaDyfcoRhu0Grf/LP
HLppMZdWnNft7Ylb15G3Ir+8vkWHK8S/pO0UJcBZUl76U8UP6kxOwNx0L+AmGVULVhCQ/tXBo5TB
isx3XmGmAnOb0u/IZ0OUt2RyOUrcKJIq6KpNkudBqolzC8amTFyWcn5o7L2IqZjQiLm+WPTYgOrO
Ce8F8zG+wJr8GXvrDUh6nWQz6UlW1T+pxky4MD8wWIoeVngPsUrAMbKPRMdUFni4u/tbifSrBFfD
h2Vx/EGS3d1015ySG5cuAyV7bpqd/D/hKbXNLDmyFvDCy3Zg/zQSai+XiOS+/vPiBYLuolXpSoV2
kAPSiYaBfUZXe+aF654ozhkLwTdxfcsQJlZKdzvnreAPSDfKua14NOC+aTuGOu0ONbEw+3JWzyKU
sborl3u9EXpDZqnXgswk55RcL0jCUWw4s29TLo9UFh2KnywlZVr6c1vr2UuUwPPOZRhFXDDXejco
7KndqR7M86ohrjZDWrVCHUo6Tot//+nYJfh07D6CsH6ky5LX9HhWwsrYHVKln+I0a86OlDaqaraL
pR4ZiNpv1be8HiDPINlwxpfadEQm6iivV/JjeQv6crYKS+rirBapPz8PDDLV0Dl28ydyKIW2g9iM
JBrfIrrH9FQPOwS4ZmDMZa78pUTHHOUOAkZ6ejGLwwpg99d/ZT0Gh+QSduACMN2X0bNmxSanDd4c
9Nqhe9k5xzEDGezl2YArhWGdDPFdy1qmps3mZU2geb2oo4lLvmtpXZv4IK8dMZvmTxBZ68BPFwBc
tnNPTZ3tqGlKKOBpR+14Ksuu2I7hb+UBWiYKzBdTBGqwyH34cOYgbKq/8AJ3maJJVsAOD6wZ9ijO
Sz2UfP9kUeP/9MPtQuPoZSTOGo3spH1FB32F+e5D2L15SYRhZjkf69+Tk5rvLxzkKXIWakdM9aD1
bW6ARYMf5GWVMsxKz8qhRm6LfQ7N2VuzKx/SkhIRlmZjqdYjHkU34E6hgTgWSLnAQ8Uue1mL62rA
h5DzbQBuYtdyxAO7ntOXrdMDguvq2I1K09U7H0cHJK3OT2g2+9qH3QA4piWc6q+EuqTnAEEQ2mYf
76RIzy0cv7ae1AqQ0qopu0dwHyw4NY/W3NImU5d07KRqCYQ3O6eWULCWUukLhHgCbi6wxOyLhKfl
B8L5vVXfjVlkZsi9XwZBh3l2kj8v3HiWerEGxZ4MLYzFokWQwzlDciTDuAykpAluc9e52XORTqPw
OUy1ZHsPcQAQXhNF1qlwlV3al3LYFIGeVtVQjRRod3QwbGF4Hl9evrdJ+36jGGuStKGZ/wtPz/Qy
Q3jIKIOYBzhzV1iTxbrsppUoIhV1DhemySWobzSGtvfdlYxxlkioHdR3FB5Nkcq72ysVEMi+C83F
G3Ol6rxekDDSFpAiEOqNYh1/fnmLhZ+bzI8Vm58q5MtLqC5qJAXdp68fSgp21dS1UlDpOCK3rtHn
/+D7GYFRXQbW3oxx06cfqP3yC+hX3kBFSbhuwMnIvyIe4KIvEghVjvKQJX80/tndcufCxPezsFhx
xJO3Noe3BsDEZRiyPAuQC+t47Y+/g/NK7rCLDlxuUCgOpdD9Wm1RCrjD7fecWGebJWdUsk9ZkuiP
i0xo1Udg/vX5/lxGxDTkhMFf9yYOQpbtoVzmHN5Z6HMrPMzrbVu+vxt6es7v3YPxY2MMrI7dMRBX
IoJ2xYB/pK3B8yFuqtsR5BzbAYkb+WU8B+fWPur4WZ2v+okFi6+1xwUBK8isq6Y8ov8AqvzibaDk
4za9QW2iXbxtLlLKZSwtJvW32B13Wh3L1lQ3SDPyanWtpNBU36PSO0CyAIB7AWB2TefSs3Bn65pO
AqkJjU/Jf/gF0aVtLWHEiwXDzwAjFBZ2C3mysnPchhry1ZZs83wOqO5+Ze+MxExVcCuLFXL1Zf8i
DdoizxslSq8Rzs24JR/NUpRjvDdqTtV45mKHIvDZ71NPCiFhnCXX7j0xGD7znjpdBkGQ/0xScPgC
ojbsYcH1E2b6qPfwbdn/WAIAEiMyMsonpGpigTYNIh93rzgXWjf3FpA/qx6AcWYigemLtQ/V5/89
AcvQDwur0yIUaLpU9xCBNVXjO6y46NZdXfwxhFij7HIe+C8G77T0t4xndn3hVjywzfDg6zbrE2jE
Xeiq8IHUuGndZI6fc5SxQDFkyZeT20P2B3OsURHiq6yha6Up744cFnuSwuuxaqRZFX4Hy9xNn9NF
mywqw368uWCgR92vL75pfbmE20EJYpDi4CWJUKCyPhuChgD21C1j8h3oA87Hv2QWOvlEghek1toK
D2At9pSu/PC8Wb6TspEdhR72Aen0/eltIbXT7/kp1QFM5kA7BcAVn7v3nbuzq9WWakpT1D79H2kx
Sh/+O6Utikh4Oy7Wc+F6EX/+mObBJxVYCvRgx/gT2GRE7157T9spTYKswHgsL3CrJGEpZH538s3j
2gEbBmLadAkEqhWuPAUE497huTrjhNQG4f5bxBEpfv5fa0lm6rZMfgVkrZSzzDSLc5rJfngUwuNB
SjV0+TmpZjOU3swGSdmYnyDTOQD7Ld3GyhYwBSR3haAA6ekkDLVv3ckynRDM/jaga3DnllthkG5I
29eTAFbJuuhcQlZe2ivF6B2yoOm05zpbFA6u2s7RHYiLkQEZxk4x9UbbYJDHv1LWAaXJXYmD53BM
Hf1IlKvTV6c4KQ1JHEDW/A8/27vpziySN0IQWLimfVn8Q+KOZWbGc4F2ayo87CZM9PUafEIk66WI
UC1qwN23Cu33n2WQXLKHZQFHkMGTNBeBuNKtNw3qdzl8Mt2HHWsD/7LlY0KBnhC2Nfi7knkD0YhV
/F+6KRjBt1S/BtNV+HT0IN7frM1KCfIFSZwjFUG6+t5DQUKBlarkxhtiEW3YyOgeNlu4vy/K+OJP
ihCE+cXRNWaCyRAsw2wUXcjMo7UaQfBZ5GPWFJKgUN0PyE2Wq6odCpQr9J4MYaB7d7PzdLQ7HTBv
Bj2OGHJTRqNJuvLYGWQTj1L+52HgLzLq/acOgv/ezORwBR0SjZa7MSShi3AeIFj6iJ8jTkhA24WZ
UFcgNQwfXN5BZbS/2Wz2aBu+G/yOK7vnXX9tn3N4E3sLTpeMKBThlzCjosYdHq3zS+DE+yB7DZuz
luOM/CJEDftvvQ64n3cDED67zd6hd5hO0zP3AmqUvnhViUYW6scwJqzIjIQ7cWSaOINPSzGvm0Q5
rbj5EkmRaUdi80A4TwJs48ww/5Co5Cyu1k8/dn8vM+ag+1dARthuPHNM8sq+etuPANvKLcIYJFXV
L8sYzQODf+sqF6W2Ls8ZvoKJxipw50yxvbr8AW9VoJN3ac1Z1D7cPfebj4S+ZHbk5eXASvNQ0i/B
aD8vZBCJQcZD3CTNiwazl+jFXsUcpd7Mgk/xSJklv5S8olrDTXa2/n/sIWzdB7kMHcyAFR0/vWPr
WUBgnO8xK55pzqW9apUtURc453c+gNRbxAy4hM/LNuMDveSGFiY7Pdm+o4KAyt/Na7BO4wYmnX9a
JvgwNfm0rMyDd++i7DvfsvNGdLX8vY+U2UZE0AWu9bqqAiPbrsuUAQngdrCvx4xNo+mfYAjMn2dJ
DC7piL4gN5uhgNnCG1wXXxGm4JG1koAiOo4bNdYGJf74ZE4AogPIGVX/VODy57BVYIra1zWZD1pZ
FvmF0GBtHa+4g5fYbwIo6VOlK4k9WctmO1fYB8+CKO6h5/oNnxN74+WqS3zFt5dNbAeW1PW4VIYI
Klbci48bfbs52H5sKBedcfsTKI6t4tRZ2/eLdxeKqu979ABOzgP6FCehk4dESLOdJTCVKKYcTZPm
IXoHtmmQ8KGosbNU2b6aGjxg0ALuaUc6REqmtgdPoH2ey9wiPYh/digqBncarXuGgt46OK54lnGL
MYmd+aMx7vEivcqk8vHeFZyn8w/kmGudg0b5+xJm/tgk4gJAaF9jmPfFLTPvA7kjdATC9Mn+0Kx8
FAIExevfvpHJq8hGxZMpO4oH/lcH2uFUx3BAV/5pv5ODDQJ63fzxj09Lm8cRI+E6T6BCqN1yiCUZ
DKygLCLdLQ8EUJiMHD2cddeiL7vNP4n5BOz9QhzzC38tsiKCMrepc7aF+9jhrh6ufqgdg/JuwHMZ
UOVOrvVbbWVToZdcaFaJZNcNAEv2dFoWrK+fqnzlOFZIL6QPe2UpKGh4GJtxvUZhXYEDiK0zIMQH
sKD6ntSBVKUM1Ihlypi5vfYGd/IocWO6EzWVkXXdcHTQ9pYoxZWejbsn7IT6cdxYU8R1il6sOeDh
w8I6w/0xPBhxB6mnMJXbTMwM2vwrv9hs6QJhJKURGv3+uXCEwSNLVf9h/G/ql+j6jINtwwdcRPCc
3isdyFssxXYMBHM7g4dfoCi2cAGhppfRZ31rblka1qblAJnDW58NJzjyNcvEiPOiPRIoyrbaeSQT
tkGovgCf9vEgSB0X2DvWJsBvokhftOTBvnybtjM9OrX8vZXkcL0RRnnFv94OxZs1R+WZTHMejleb
x1ugJrbtRiAG8lCHQ1z8sLpJhrOaedEh6hhPYLNVjh/W0rrer1fTdzidGyDZYSLSOpXOCouaBlu8
ANCp98xoluBgl25H1Vt4U+cuK4SLuZN8UEItjtnr4wh48Inx4Ut9tlW92NMM5B1zIvgmvWID+fF8
M68mblUCS0xB9eOREcIbE/Q/+aIFz28eP50h5z9CwjO/Wlb8aK2WEtasOCrwTxWdZDTrm4MFN36i
duRV2IIVFtSG78E0tElzfpH0DgUXG0VGiFIDbXCSfL8Uaiy3Wgy4GNexdPiRZmW+EipEMAbVG0q1
fRrJW1sTPWX+/5iJuIy3zi1+CyiiPtH740P3I2kPPLvInCi/LbKEIgfuHxWS3LOSwzTRlCCBq9o8
DzvIaPhJfRPPOeIKYxDcXyK7sqFl1PEYWYa7pFMtxP+lLj2/FqDd09LsAgKWXs1pDb9qrgk1FbqH
PPYC2ppM9tlHp7WiicGv9c5vOTuEXV/9AA/4KmJuRPUac0RD8EfFuBTP4CgVHrZTOAHh+yH57cdF
Vc3EiRz+k0rJh/nejhZFFPqhSGsLJSCFlqNqTNue4txrJSVAQXIaugmcpGyeah2VEOGPV/OuqZGr
n/+WIxIWtpiYMCoePYtLljJpmkPI5AwnyPA5qKxiqMxmfoKIHaaKldJ1E9duMJyhF0ocli70HvGv
bXvSxCUZz14Q5SRWySMWrs/maX2PqqEEOQQJcqiWD10Zirk6Ww11Qrm5nK2Kl2qzY7SEth120V0g
+CtlHmyYaB8MpZaoGGVSoMnMLsp1QYp1dViDNbKbYDMb0c7y6r5GQTs4NGpdmSN6BUQvytv/ELCc
+wwm0ByV/15ms2xcyYejyIJUvHZn8alSgGsKRXX0CxscQqI1IT1XRcOHxjjJOypGhcT2NH8TdzoI
9qEk5oXpzB+fT3RkwmfRmmWC+jj6+2g4ySQR2OXmnA35RXdMxIsNFouUGar9xaCjsgftj++Kv6NM
k+E0DzzohPwa1nkU0ROnT53VqVYLnaGv9fTI49GZ+mSi84JW9wb/HoYPoNeohUTiGDYSIhv0EDo5
mLH4h/ecF3t7FoOKEY3wLSqrM0oZvUtA8+2ovj1VHzBg1pdP0NLYwdOdhkqDErguM9qupbv6TBiP
bKYiOjVkhU1MipnXp4pH3tl6KSjzk88BtBi24Obu3ZB32pxP/JGTJl8G9xhDiwBpQcFfm/mpHhRf
Ai/jAj+3wjiOog6NapKAP9bB3l12auKGeb3R9RFr5WoK14KYONcc2me0ydjsUXecbCZKdd2gL0aw
IyXInesy0LRS9EWYAR7dbrMFltCssNwQeOH2f0ZQaWlWezwrDTPSaqbBn2fjEDr2GFf9ZNQj1FH0
FNhUjnczoskiI2EVbxBbbkFLqYMjCWbdyn1Ro6aaBNzXRDwef2adxVOneQN2w3jwrmlIifTeKqgP
bYsB/umrCQkwsu90gbiX/kOF7xH4bJyTyjb9xFcO35wfO8Xw9mnbdTULPtEWvsDv4+oqVOAyfwhq
Vo69CM/peYVp+Kgia4MY04QYr2uQ9HoesbI5sFtBt8v4+db6Ht45jTaiSW4LkL6izgjVRur/gkK6
BjwjaCgAVUir0HeqZlZkGpxGf7yGwo9w0LsDtnqooTfhcUaZgWNhZaBhDqnLjDNcMZ5G1RP6Lunx
0FfnPs8fgG9yrrqNNZNhImSNry/5HekMmh6xgHru1bvSwbyFcaEPZDzUvQXZZkyOapsZ66UTI47P
Kw6HsZn/4DDCOomzREyijn78oY3uRx3mJ2C5X41Omr9G9eNS3v1GHdXuSDWch03t/Z7D0ma7sfnt
crmuye4LoPFTGUsSaKrO2WX5rftmCv0k0Ht4Ct5tiwDGqdaEnw8KlEh5GtShhKCO8Fg+/PL6TAgC
BKxMH4Q6ZySSer9lI1BbEZ3My3WOxf+XbYTN2tkPSGJhWes8k1o5K0baFf0PpHD00OL6oGRD/42h
IEYhxmjkY/yAAxIk464AVetXDCUctAZm/TOV5+jJcKzj5FMFrL1Vtek75CQlmkZt+eRCfkw+xkNI
lp8d3H2A2sZETbuljG1/95qDdbEjdmWZIpcaF9yMMm3fSsAfNa26U5fieK8Fq8Pxppzb1L5QSkik
66vdZo1+HQcWb5Rs19TnGtLZt6QZl30lnbuCFsYmT12TrbDXuy48LKpeaMtFlSv1Z2xAPpUSju9I
LuGNn65IWA+EDwo+5CfG+f5S06AI0BChfT0P0XB6LarSzTGTiBHbOINZa8X4FT68yhGsLTbd86xR
V8HlSzPbPh40owyA/5U6ubKh4T9dv0d1SZR+M5dXqvZlLGEX0o/6fXjueBrrrXgLrKok9aaika81
x5PClVwW0AYe5HkW3FT6k5A7s2YGaJBsVQWseBU/u5eyOIiw56bLSPNkkxbepMQPfENWTxxWE8I1
DcJT6UUzrlZQQchfQcfHyUJ8tw40rVOoay8x8fe7H/31/dalbJfVBX85Ba/2P6a+Vul1pZMkoN+X
cuvPMP+J4A4+9LsIJCp/VuOBM8o5SluX6PFeQPuAD7xtUxL3h7nmCF0e3Og1EykTZY1LaQBTv/BE
IRN2+ny4dcmJz7L8G0DzWMbRbfwqy3ODW2a1uoYumgPT5MAVUQqcu+O7B6Rt5lSrFHyVznsueXzv
qBrnjCCWNCO2XoZwcsflvfUOh41oy9wm2qZutLDb9ob/TlllTZp+NH7H2dBoM1Llj8wVR5lL8mQQ
GVGgN6y8oLCu+ccNjST5NIS8JAStGdnY6TZe9xUD45CwkhsJ21m6FIzPEC7hiDtmwdGn97dAkYkB
6IC6S18CFXqvNrQKJ4sVrDg8a4Wx8a2U9v6K5OXs7MLNvDqDdwyp6LLQ1GIutDn9LvN1vOcOwzwr
pZtTC9eXXGTN+hPCfQ7d54JePUFXcwUBdoyCghrrzOVEzOjXzriaiPxEywVGZ7pKEJ8LbItDt7jY
45e4iAJhIe6HKUqpWh6m6+Kxy/Du7DJ6RsJVnGb+9H2Tq/2N1tSlX0Tq84sOl1fV/Sv/yT+ip+IX
gD4tABv5teQipY2VPIddp7TmcYGGbsAYcSegiaVVeghqe05je2r1XChJlfukW1fAqOSIuMBf8EvO
4mGO9bsOcx0pNEWG3eN3HM/u1A8GjTSvFKEmqHDTEhIQ8IvpWzvkHfXsUAgueZi3YB+ah2ZxtfQm
mqkqg5qrf6af3NpGSvU9eUv+yHO0YN1TT1jnjaC5yfdRNe9nNGVnESNknwQ4zCyBVQGkfNEP6rKd
nkO8Gbjif2+miFvGM1XcOIV1KgsJxqPSHc1CTl/3VSZ40rXn7DnoIFgI80gSl0cj/LyVpoJSPF2V
cGLLffzVXoZn2+zfR1dHvC6eEpqF6b6+rtTbFwbKZJyKMGKTrvf1MFHSYj/rMsIx/3g45BTMlg56
6vN3JzJwop0XZZiKwDxYLFO294xaJnEpU7D24MBa906vzTpDXi1XlhT8IJB/hQzdzd86ZH+o4NzR
8Ly4dmryzEVE0lX7W1LDs6jHYRmfpor1yZaqJoTL4RtCPthRbfRYwAXbYrz+3tB6PJUI1jXr57Ec
za3IQXPloGcA8EuZEwcGyCCJXnQyD1y0TCWz3gPSeWRTB03xe7juqvxMnpgkoDEHPvU4aYN/AxTh
RDJ2PyFEoCZMWYY3PSEW2IpXKPx37uuW+7GWpht4Oq86qHAsWxtlsJ+lzHRoF1RwCc3+HjjtHdvf
7oniLtNkNR5ueEx8s3h9wpLlG1uPE50j8Xm+tDUscqCpJXZ/FPimWCM9Khkv7isHghbAShKwDjx+
PVGvY3Eq7d7GH1Ge78+tXLWUNKd+fKH3K6snGTBNxQ4CpAkWRPZOPFEfm/6l/9nlLwbeTf1wp6vp
QKS1JCQxUva6rtaeLyLEnH2EPPWuLAxDVfUtR6WtTItUYu2YwrGeAw376po07f1nZLPoA5KZ0pR2
WoPv6Grs3iEtDud/h5Gdj775gpzd38K0EodCpwxBsdms/bac8SDY1g4zqpJBcWvoPEuy5pMyJf9q
dPPxUK8GqhLZ8t5M3hRHJ9KXNH/giOv4Vg5rZ8wYCOZF6QKYA5E2w4oiyctbccKu0MOhYcnOAanP
H6e4A+ayG6MGdw2Q2RZ721zmRg7cSabrG1CybRNNOcGc94LgTPiuS5UakkmF341RowrFPmePs105
bHB/fevUY6UNd6KoE6UFEAluNYU5Th4aFI+9/64vTGZOypuTnpxLAKoKDEC8Qne3NGCmwPYPYuI4
HZwXe/Z91JYTLAB5qXgKntH+yI4v9rVID1Dne3OtHjoktzeMhix4bfPtg/pdp825b8GLj20YOv/A
N8sYmIC+Xp4shLoQ4SXWjMhFEDfAlDm4FrCpHTv+YoodyCqJvuix5DqweDRz1X2c5+Vw+aK/r9bF
0YCo5+gUobKNxnpGhl+go3MJnklRiewuXJHYnOghSmQxa2Q8gLDdgRffGK7P0jy1AZiYW6JIoyoj
ltfNp3ksgNYuiL5EAU9tsn9TU7UM6xvP8Cg6SvEJrW1huCBcIShz6uATBT6vunRtt2DeNEdsFrJT
THxghL9wz3QHhQeb1iBtFRHShNRwf/06jYopHPDKrC3VHoPJ8LgEjf2YUp+uI1pHNpflMkuVcL+F
MuFuI9hSC5b4xWw6mYpWrFWSPUcIDltGW0OsEefT5mloRZIRsF3M07TGU1jnyPvtUteUQUZIaGWQ
SIGr8emZ6NZBuDyuBz7H+8kRM5DF0OThaJVA+zNxl3NsQf4HjkEqYnZ+X+m0+hkS1jedKSOJJ2uJ
0kMj3x9n06A5D412BRhZbA0TVyJuDgEhikfqXHVOfueUbwTaiR1coqTJgmpN4LPRXCJnkqMsYdwT
ZkmUT41uZfIaubhPtrlxXq4drmNbw0dZCkJ2KQEBY5tFHTdQGpYp5UdA6tLfdHMrHvbT9enYT38g
aJHf5SAzWdDphQts4wlmKZ4h2ppMOy/pxVQ1o8gYMjwbh7IU4JA4Lq1sbqkb2LsGBAELUL8JxhKs
oGfSNYE5wDC3UlktyGG8cyeNWXR/Xd+Nc3RkwWfSEYFnSQh4ygkEo0G/sVB9MIAZcYj3vskJsDK8
KsdV526NJcrhLYh68WAan0m+O4+6jbomSiatjq03mGNNnYJLGrlUnVJ6TpUPyJtqSKaAdmLw2aud
smHxpxxswEa7JMwXvlDc7AlfyJ0nOwfON3WsxpblQU5ckVKjG79m8anh/lnsZb/aCOIpHoGA9Hxg
JKUJiYLCrLLDGz43HKUBCmMft0xK2VGj7BBU+FBx9HLBzmbCtilHxffy4B7dFMHs7hlAFv1txgsm
gBpOD6bCyVhH9t8Uc9ll05NHNvzhgW2pltfcwQFYp82kzZNt25CotBo5TQ6iXw3w9wNQwbGzbkWE
cVPCc1+9xQdZbhhTz7oeFtXo144sRJBkSRtpJrEg68IWEroDtR/wRWQZs+4xIzIQhYzDoyg61j+o
miHuG9muS5HRuk+YUybdl9YBmcTAW5DLbnoyZLHqBPJBrMR6nmMkE/d5a4QkSy0N7XKKd4DylYhD
/Zh2Zp12XpqPap3oI2vfLxFctb1B/HlQ7vIyl/bU8rIGjn0BCO6bwM2B7ya/mwS+rbqddqWMQYdE
g53Ycf8BCkrrsi7UMmXeV5AJMLLV9ltxTZlmxEoK0xOSTPd+oBEkBRuauteJsKfCjDk4/vn1YQju
UHKTtQb8PjqRw7YnJHdeQJu2Rz0OeYqGrMqddbGM/FRYKqanu4IlDy9J36uFwpp1E1+iabRRQSoe
v+mKx2FIMOKs7Z3rN8KgmjoZgjWEqXlrxAb8gwwOKaGBI/F8qaHT79voqi9DXwD+Us4C8dHyJawT
RbpWCeMzDIiq6fHi7ybJFygwAuheOYoeOZZRkgEAelqh02L9oNdB6J5JQFDamK4Bmne6ukvM6qfw
HR/dnVpTPehSBupgE547jSdbdtU1C3NfMz4PUZwQqO6s0xq3s4hRABNPBunPTf2Fk0aZ2xXwgcew
okejEZCMBcobd7eii28keI0K7+pc1lGTmJ2gwtpBKkKoMB+GMhvJ7bFj3gUm56YmlovOx6NnDBRn
nibXK9w7ZcX7u9gaTsBVV/3UiJNT5WcJD+IfXMIrmannfvNjj4bfIELTKLJtapaKUj3so/eOR8jt
TkTn6zjkglubTmcewS9ZSVh3P6n5VprlsElep6uZ9ZmdOYeCDHgDexZ8Hh4XZBL828aawH6NJhY0
SSjxGAeoGZg9qN4Nr70L3JpcaMRluKWXRlKROpy6BlOIVKbIr6g6OgtHZwnYs9mtuZK9NCNiW/DJ
3iMmRV4qe6Xo9tUPaHlt1ocjVYOJz9ffmCn8faievUb8ZUc088EfXXI8FXK9o11UqGyULXMOvELM
64oMl4g/qXYnU0cv7ruN0w6Y3RiW9sxCvn5GdL5qoN1FJEvNMLFaqGsgJiT6GLzE4qpv664+qXFc
Rmol9xNlWdUCbnNGBWx6hobrBd6kWFYI+qHcUufDM42TjRRhJ7jxk41vGE/85IbvUSVcWmilQ+86
soMRrNxOGjwZw+FX1a5Sbeg3lcFMsSgVMudZsWOeyLzjYLVG0j7twAo2Jq9GSZLoVQ/qn/FmVLWc
ltu75m/+BGhjGrMiKCZm2fXcvpqerxbBvYYcTJ3H5lkeYQm8KHN8a9PInvjo72HlDPvnNKyBQHKH
WTekzEqfif+GnmJPrcFuNrZrif/hvHsdxiK+oCdJYrkNUumDNAnsOiU90EoYfL9tZ4etmAH8vUym
d2OviQXBPaOMwzx53TPbrtKHFRJnPqusbdoxcvBZaSPl+uET6znIJX3K5Tz78qG+n0/dtzFsX0wA
+ODlb69U7we0M/ARlZcTucYZmu14XX1S9uIi7hxx9R+Npzs2BC5VQXh75ZoYIyfOdkwu+1II11DV
qnIVyuJ82Q8FkkQvqRV25J4mtxnykDaBODlY1puptfmUT14nxmzsAM7nShrxoAIogERTysNRjHdE
tf9LWXYP2xDIuqmag6VuOIF1nsYarVB/Twd+78w6GFufr3EfmbSA0LkaetWgj3xCrZAugFyxMzij
o4y22YKv0BsypWHc4F9w1Z96pNZfPwUXlA4SZ4ZVkaOncral/2AMxE4X8SOXmRWu0eMoi4Q9FUQo
hb9VjLvU6B1qkrDvCGw9n+QPvODNuRRwhJ1OxglcnJ3kd8O5SHmQ0f4hfxaGqTEepozk/qySenXJ
24iMJIIAxg/UzxZBdl8a9n8Wn6wU6cmfqN57aaCXUZqxJIOaLJN1EvobKcw5krwtUZwrAF3sc/Kv
86Sg3blVPfiIH/yS/kw1C1Tis5pR1Q6RWZZtQREBUAavy6M6uFOgKKsv2HfD2kDZn8xAbxPHdM/n
yo/3bNW0rUqwhlgbUoscdQG7Iael5FHL7yi/aZGfj0gIWp04omScyPhloz+GgwCMS0fG8HQI0itR
6PJtnPk064Mb0RelbANZF6oSbjpeV0EMjOoKPRY2uDKsrTVoi4ohpIRkxvWbWVFmaO2EPTfPQvuK
vtuOQcwuse8IQwmTeV2GR/0noXv5J3AUEQZgDgBRoUUqtbSYk41Mx2HpP/nuNVr6a2OaDoxmL3vb
A11HMpSWr1edop9kpp+xwrF0UHnBm2L2iFMJK1wB2/CS7mSEe16JTEu0NsyF1/oojRQ+K55HTiLT
8t5pW5Q4tCfwcsPVxfO+YtfzUQ8UxlvdeRJp4WKb4idQHYkz8SwMGkSpN8E8ETwJ8UDQm2eph6qn
o4+AUA1LN8gXu4Wx45AIdTpGruV2oFFJPkkMQhJXjEfBmbiL619jNn75Pj+ZD2NNgs/6QgJWV5a9
kYL7OfPTaFdiOvu8OcCpEUMsCZR8Nn+R/f9M3h4TEWVew/d5eHzyiD+Oh7cGVyGnZsmfN5W5jV+l
0gT0feyu+8ej/bi7eRLF4oYkG0eC3LSVXZqOZu1viMqA6rfqC6tOH/xUyXmPYclL+YFtbfrIf0uP
wTWBtYQOX+jWGuFE7Mx1bAxLE9+5/70y2cTFkt6k59Xbex4jqme/MWx11+U1pK2UP0dxP1CWwMPn
WDoqZs4MnyDC/riLah6U/NJsPwvHyQ/1/gYeYjBAXV68cEnuJcbh4+J50IBK6PJWILgkyw2S/waf
sfQRCV7JHjFP1HvWveoUccXGr7F4CZBoKW61aRWUTl2bZ4Z902JGUk6ih1vnBteJ5Nh/ljigrzrM
7oEEODQDuxqiQCezExI2aYn3a9qJMEStb0BYz7rVlSxSIkuW7jwInRRYTu//D3FKga3kIZmjX/Ur
UKLH2Fs/xbYkJjOaS4qzfxUZHElN8ZYhurNceippVv0KvZwEWvBfdb6aTEqZ4jbzk4r+gX9ANHch
5ZNo9cbFxAI4xc5PO1eF9M/4MIdafiOb0wFBNFnxu6fN34RFzbYJqDuZ/O8CqlH3jQ2u4Zht7/Ej
wR/1vguR6mtO6QgIaqeGd+Tab3/IhHk7CzPuqFgthOlZEAFHt7wIba0P9kQTOIVGtAJw8Ylto2nP
RCjQSqxOqjO9pOStABtpVSGIv6NlENSyQNlgpaKElSHlmrP3lxdgGJuPpDxPTM3z7cKDzJWP38cI
JhfzenR4Rg91jMOzTi6LTFoJSfTjAF+B2pfrMXMMUz8VsOQ7dTFyDIKNjB8i+NHTh2TN2umYRFaw
6ksXwc+hXbVWorsn6J3VPjb8ZE9Uw8TEsO7DvqcVGBV+lvSNzgCo9dyJZE6ybjoiESESToxNmxGO
G5Bdr3yQfe+PppB9q07GLXjCOenlwK3l9GcxcgY6Dym9/wx/umNvw66YMGdm2X5zQYx89rlP8R4f
Rk2hNKbKMkBfhpi3iIuaSQZ1yRGD125c4PX/y/1k3V/P4sBsD09fT/HLKYUZwS33cOuMg/nSU3by
YBMHORG0YSzr+93bLU+xyfimuAzOYM5+9Jq1eAWDbgVBUdp7DPWbqBt+uNtn2hr2QWuIi/ekAoU9
xyTFDJhSm7k6vMZnpenB6SdPSpMyKyWZM4PrjWblH9gOhARdippp3Q0rQdF2mL3rsvSi4Qt6gTA3
nM8RW3pmFBF3dBTZjg7rx8fkvFl8fxkr+XPYIwCpFNDSac8ThQnGqdvDIPKc6jTpCEr/0whkvWyy
lLTz2MbGqLRLnNWuY2MGPAtJr4EHZCGY1YauxqG/O3KH9ZnW0onqDZrIGtYfvKq9dFuUHXGg7iAR
afuiJvCHup8Vc/cmMMvBI8a0X2vq9T/6RLfRARy9+dN5ahmagetFaqNhHQ8rGgrgmwZ3b3AmwxVd
eg/Ulva8aVRGpDzcNIIG+RgeF7GBf/5SXXrqE8Zwnkxw4Rk6+vq9X9oaJDXy4U1RSmV8w6W2kUS3
HdkV4X1zmSJ3guViEIzCbpwHiH7n8mwM5ZW/ddhAPcfDrPuTvFBfOjULg8GT6E6N1vn/5FjuCHq3
OPYs5xfoObNEy6nAlELjGwaAQPLzQGkAWtv2PDG8gcBfAh9R/vfzAhOrjVkYKEqHogd3wEn2SV5z
OBDYQyWp0KmbGOnQeYKAXsXm6cfBIZ5MoJIfE+iHJz1j3+cq0/7hzNQ3nyYmN7c1GRmKn0dmREX3
/mWWVUYvFwd9d+usUTDvErGv2L4e8G9pvS20zj4jn7MnJuGCDrn0le5o950pYrJJ3SzuMG3DP387
q7nxvYofwJw4xlLJQ4rZ8zUpoI/lTetK7FUlp6eaku8K8ItYIO+ppdvFO02Q5FC3e7DyJ5Rv46Jx
HRzT2mjX+D9VdHNvIbWX7hEUQ193DmHgVJt3k8L81MVhZ4EUGfk+vTgRuCS8O28Wzq/cayfqxADk
DVOPymUscVATojkB+YJw9TzCP9/fyholGTp4Gnu5CsFMLAdWP7a+HGxjGl4vNyh6s8zt/sfmSsvS
LOHu7GTcaZKdXnzH7gwVYvDMGi3SiNJI/O9hj/sRwuHLcKWKQXOBwdE/jeypVkB0MMPhxxFToKFY
suM/839koT94BS4ZBuOSV79W90ZSMUlIPSKL7z96dlKGLfXrIN87/c0yItCz5PSjMx3YePyq19Jh
4LRLzJFE+qa9bydaqr0YwDC+ftIgrjjJD7tdEN3cUhCrm8KgeoaZTT0n3uF0oj0EyNDhDReZ/Rcg
iIlxIbwUJm41HrhIGNRA0oKnb7ZwM7DCDM4oRWq0nflqNoTEwEYG4c5YmbgMmQHHDVW1KrBmweu3
lhmwCARpx72JmrQY337Iv+xP0CGOUoum+7R3z8WPGpIDF6tzH9TgiEgHMJRcpe6jNwm+Q4ipOuaE
BYsv1eFoY7vmiLDHVcUyiCaeRYDfUVtp4LfzEakgROAPjS5JFzMJ2w7S0k0/2UsXhKeQMInM2Mv1
wFuR73/1flrPIIhWEzBuS0v+D0Fub0BsuCHwLjYp0rYoD84bydaHfm8Zj6trQKdBi/hPls+X/yND
NOzKVd2SvpAqKHu4wf7JGDmGYtkzPIwctYyq3lzzeIeAW0z/IHQEltZ3yxcvcJ8a8bYwejwUoUpV
cqDOBMOO3BLWCFUPqcR9VxYhM+bScYjyJwST6pfSf8aPcxcUWjJuoY/u2+No9iM8p7at/dIGcjEa
6yCNqyCCjdZMgJ7CNijQYsCzj0Us2vMp8ukcrIXy4uPA58dnQHYXiHDxGAkC/d8QKFlx29nsyKqt
6936QQlo89fyF5KUlUX09VRYJsFGvbxgZBGW2KBhH1ARK96J4N95v/sItYzuaghxSmwI7FUkUZYk
AVZojHDzB0OZvnTrjb7EUuIXo8SNnVOUlhm33N/osyVF5NDOu+ILaR7Xr1XQTmDh5Pdq3Ycma4zu
esSVpRIyBMBv/BLrDcMP6hdnulHJns5YS/B/lfQJPS6kSMbt8KXO0QJ+uaSmit/LdxINJVSTTo/P
PTKfOlL3InoXA34v5sYWTze/fj0HBtBjPYfIc8laEVOMhx8kA5Z7e7HJGVnou0Eb0jBbJ5pxIdJv
Tnc2I/lVBRJE54+W/L+sySHVC5euTmDcQ4f35I4xePrvXfiD1Mn8Mebo+XXNVJm33yxWRskJIfcb
68velKoPqxvXbj2Q9G0JDzVwZINXmAVsNP/N5nJ+z50J4umyU/z4dHBrEHX53QWey1ZFtdVHTogA
pKf67KBfzyPuwG+HcZfK8f5E4ho1s3TafqeqgJR7C8QoXkxdRYjLxzk9mU9itwdO0jrrMamBFB+n
PRkZiaQwm4UahljCvS1eDiXVYKgk610zWRjM00jQFf0+1GoJ9siDEoqm1HyoPKQwJic6aX0lRqYj
Pl++tBURrVrm4x2cT9rtKB/g4k1hgxV2GvG7I0GEqhw6WlIVPdLswHMIqY1Wzygq+O9ZrbRCHS8s
aQOtmUBp1p+0S+0cF2H47WUW0Q0EmDx7ckly96Z8NXkik00KnqWS3vZcPpVdhJ3aiUe8Jsl/7lSq
olLv7DX3FVtH6z4RfZctef78LLeiHm2bnVbFrIhdE9qHGRC9DT78LekIlZPPWijf+n/ocKIvbGzw
8NxWxgejEKAZ69MdVaNK8WethWwpt48952DdJ1JZsTo7T3G5cWfSvDf65tBJye2/sYcq5moAfdAb
5LcZh2Pu4OMyKan2pPwxTXGhOeIc2A5dWY0fN9bgblTTuTbByuzFTjGaAofsePNKw7AqvKjDt2g+
nDwUBv3g3oFjNliy+bR3Dv35Vmk81bkFs7VJ/Lxvyuj0/6iVB3re+Ecwtiw5UIuvTmsVPEQ+Hk41
+ZYradUgubaXoeWsl4DLjhILlGBZyS01YvaHlffCz8c51xmIEBo0w9gw+S/0ondX+DTLgKiVAlDS
ISJZJ840aAb7XxeKa9WCFtQ96ZbzSYqhZSnmX5i3QM560659o21+3SBzCqrWlNhQX4+Nh/P6lQaa
JCSI6D3wt1jfE6YQuynESfLK1x7TvQHtws41Grsudz4obH4WKR3J+xYTrigTejmLpLOAzdVfeMZK
3gfUNJpDaZSn+wnkIeJe+K8D1fz7yeyAyg6peoC+QU7F6tWdCizMRX1yiLl3uAiQbfSVDis4lVGU
H9N42oqkC2qAaO5goX0Wd9Ce/OxGSU6da/e5y7Ui5tDyX5JvzB2Wy2Ub5WHeEymModVSg/C7yXi+
ykDeB4Uofesf6g4wYemKpgXCwNp3426KbFtUKoiHAywYJifB4QibdPu2YIg3lgCMIybwoGvRFrTi
38PrjgETtkkJFWkJuAPL9CPQy1FXGJypoNnTLKiGVTVXSGmIxMMIbn3oOZTvd80rlMJeXgzTqpsZ
1t64Luxq2RevQvGql5Glg7lnTJpkFtLK4SK0JkN+Jr3HShueIq896goGtKlC+LNHrvID4uO5GqDb
2X4LbPOk/el9u0p2kZ+1BfIPArDQMaDXzETp1QQfoII0Z11NoOu9lnTsPDe7jX4oq4veOqvPQ7tI
6TpXusPqWtvcayO5H2yWuYPcqneLFWra+Fqix8+8ai9629xqUCoUQjc865gji684h0R7zWHJx4EK
xES3koc+qAhub30rtf+GDgsG5YlVYxe5f+oHWeEKkl2t/1aqkif/v0h4kr1Fv7O0GsfxcmxM+OCI
W4JgOFlz8mUcDAqhqn54Qljf0I6lukwMxYxeiVBp/fOD373IICDtAJFtMeeDOmPcNrUCo/fOTuIl
gAtzbJZmH76zHMRcznpvhVTTHUCejKKdH9/ec1/+ZMKn9kyvsAcE8GRJud4Awj4GyIkDLWNqCgsS
QPYZt28qcCamxpxtD6WeT3zkWSTSLluJtAn3wJdyNnBhOwiuku/dRO9JGwWLCVxC3yNKUssJjGef
6awiXk6bYucDVJnV9uRnMBSi4Jv7kT0yNdpRZTqLFax2Bf4/P7EcYFP9wKV79ibRcehaXJlQdnQ8
2JHnsKSciy1dMmIqmVHUBhqLnq5qv2exgAEzEqaM8on/PXxOaG4ZqxIn2XwdWZWRDmnva9t+E5C3
IgcaYAnNze586PrgdUKuwAnOnzieaVJYnpo4c/7yLrFA2H0Y2pVZJlK3YskGUdGjTccnRf9UwjPX
YsSPgT+lMiToAA23+1hAMXOEQAqrmkjJpwyqepTLoZxUDP1H0LRKjYvLX7dq2Pyufgq5tbvcOQeG
BhpDFZimicNS+12arWXqG9nFyvdQ+nwQt2gZXkLlgpvHSa2yhOTJqMQcdqFXkb5WiYEmZKGG85bl
9KnHO0gsRFrFjJG1xfSqnWYgARXP4DHgi0E+mDIHgpOU38WvpH3aUitWOgrzZMoDvBYRScwlfKsQ
i1FDFaq8kluKVRWnYsvZve32fkx+bAou33aA+sXZdZLSiaRu2KuzYwnoHv7YTOpd/Z+eIKtorXtG
dGwKSDrHkZ26g8OPWq4VycO9yZ8FiMHfEaWCcnx/vjX7SlGAxNaSliSp58L6v0sVScNSEzFr89Fz
rHOAIQM4QjnRqkr4tMm6Us+TxLVpOSOu0VeeHk8nrjKDZBGIImqd8cxJWNWhArIdWFV3UG+fqfWU
D0+QqXbsPimBJTkQW3jLs+TlzyusCZ/UzH4qY20QaHw+4ruH1kdIK6y2GFO2Lqbie/2LQ3f0L+17
/f4ltIaoeK5kd3GeDfxuhz4trCZCBZAmmAIlqjfMkgm7xLiEwyxVzCo4I+GrPgbIy0/y9l+fJ7xA
+s0vp1ZQjiGK3cj3MLHh683ihV/9sOGiyoFDAkOIvuRrKiO44X0yEyT/JF94pKRdAiBJqgErHFgK
ycU4s9LaG9iHk/GwpkqDucMUrqigYsfgOAGy3dWIQ12QEoGXRqdUcvlnq9H5Pm2tdCeAL6tlJOGb
SyKlc+5A2GS+A7QUKnDiWR7fJXLIvy/XrD/Bw1wgH5PB8puRHhsj73mKkXJMDlFT0Cfg5gaQt3Pl
pxN/I/hDOujwFUK5ZkeuNEJr8bWPib7dsGi7ms+9M+5anGDd7AhtEXL6sghABslben/hjCHuBgkM
PV3wEYlHQ1GJZkTjFBcho6qPLXo/lMU5IoanT8mdFUvrLV9W02cQUYy0q3ablq3sY0V0gsU0TIo8
HmL7B7LnJFrvWjY8VISNi1e3pPxx+NKFpq0oMKuEUukZKhMeV1uwgG+PTPvc8QFYCRjOYZAirOLU
ZsrOzVDtHVmVoIqis3+1rXon4njWInhQptN4+37pdyori8qmOcRwUL/lPtju9EcI4EsjV/KQPzLe
Kzxa+5EqA5cetchTe8vcO8RvR28pIvASe8qnD+PK27nnYpU4DWCVNckRGvBXJRw5xYK6ONNiD4Lb
6NGJQVl4NeY4MItLZ9b038elY0rIMoZhrUk7ULWb/zCaq9qTCRH8fWtngwRHW1QDfzpt11kJczk7
O2n+Hr/czSMQY7Ig1nYWQwxSFhYaQlORo9LWr/iP88pemgCVikMub0Ncd/nVQr3WMJbH/qpFArWn
rEbb/bMePrAohBNoSGL9k2WywdwD4bFNbrf3y7wYkaIPIyBLWj/DCGaNgtqOgXDlCn56QItDfFrO
5BZ1RBbGORTaqdyxsdkUWnhcdjuYWD0cx+vx5T9cuCB6hlb05GgiTzkNsjQCy1Upd6NhCLcsbOVn
XOVoN1SeS13snu6KVIXrCVpNOiBCdWpXvAGls3csbCYJwEJW3AdKzW/w56JFNDMI1PkDfoEE7K11
qu2Jr0tFN5l8/6SffP2fHF6M78HRTMBSR0VJml2tcUz5Qxu9/OTcfmX0DibeCfi7d8iZkE6cEjVQ
gx1ItQP0YZuUM/ZQqvkahs8pzrDJXtU2kFMy1eANfS3juLYv8Hu9prebJBorb82yDrLNamqLYsq6
qDSkUxDCrdW8Vejvf2A8BtHLu5TU0U4DQp2ZP4irLorl9x+4b7P2hj92ZAC5zyJS2U+fPfLDA0Xn
SoOJyYLJLaUjKwPsfDwcT6Q0tTIy00ClGyEo3VnRfa1J+DIoueCPV+tom/4R8rdHISBsMENQUD2w
mzarj1Q+GwkTg2QBlOaks5YLidPktMQS7m05cbL2e0mDfk5Gm3+7Qflaau5ORc6bs+UHY/1k/Vv1
5p/n61tMpr195SrL8B7ZVQJ1C6x+IcVIC9j6rNoQ3QgQN4AsnDNn1pVTaVDaXvnmnJeGzgpLuJaO
RgdYG7S3jgjQ/XV2H1Mp/Yv1yOfWjd17ywFSMH0ek+clouNoum/UHEYt3m/jliWIybtikzxfnwZq
fJpJLPl5jj/NNU5CXuggnN+vSRzqXJnFeter3w+MPxS3ojtWQIPf5mwTjYJzE+4tSRI9iw75OYBo
j60iF0hULBB2kbDqRCKTxW40juX2Q3T4lx0Vhk93W+XdN7RBIsMzQJhP7AqAJMhHifzGat5LAgcN
WoKsKp2WAmdwPBgr5tHXuzNRJcrDYzbzAPAtWfblSpVh5DbnXouztrYci1d/ftj1maWssB79cqe9
A4Fi2b5YwOBCutedpXdL+ShMrtvHoVfhrTowKmrWpy+aazpf5etHMeoWQNxaTR8lOxxvTmQP14hZ
WSZTv9iR3u5Xbw9KLHKdvKOto8az4wr32GaLendFKQJLgNz4KsSbK/HVdUBJ8XQcBcfrXQMG1rX7
wTU5q2ZoUZ0O1+Bt4LjhatbIPi3w/z7QDRtEQ8a63iWXhN2Wc+v+XkZu91d2qr6knvV8bPt1N5Nj
GMfIy/C6BxJHSYeSxbd8ERPUn/D0XEHUdK/XogSFGp9Mq2DyU+ibRpE4QAQqlFoxcUBg50PuTySY
E2/4aVTD2cJ57Pb8Jy3pTo/FZYGOFqcPee51MuQ2tnOLdQwERvWwTKhMOjcc1d7i0p0Ks+MaJbpi
+tqLPHdknwBqlkBZ+UCGY8OO7aqyVexYuMoE1gCUNvPkq63wb4xv6q60afdN9I79vQRwCNUo8Bs+
4fFCbCd0gODJwpeoToOqDhA+XK2So2BubmGNznqPEwPXUrT0hFTSrhngMvhsPjPG91rSHl/IjMyQ
5JdKtvUhuh55LOuzijZ7KLPRWg+jzGuIlbUpGo+tB8gx6n/AGpt7qD4xZ5IrjeK/tw5y+ap+2ui+
eIZQhsGr+rpo+0wU7JyUOl4lx6BTLSt71TSZpvDyAFMdpd45lFmA+FUW0Ncly0yTjDwFjBrlqvKz
+7yYIGNCb9pFVXJTaK0k6+/BF1OBWP149dea8lCTUaoQ60iVkxzv1M8w6TK9I9SRdadfTcXFOGkO
nhw59rVUFCOFP+rJjskdKlUpwTdEkBBfGRx9dxlxoP8GgSdn9VzpvTFZkP+oVmC80ocTolg+Kaup
b4rSLCnqthDx60B/6X85EFAHS+i9PGiukUvrsgnvNIgVsNxzSFspIApc4ElWlLp/J0Ohvp8i8d/Q
T29JNevPn3fJYDrl5bky4TfUEyHIZYy12+0nu6P6OLljZWeOdCnXzID+/eYjyQ0JAUFR3Tzl7ix1
NwE7DbXOxheVx0/q8uqTlZIsY2eNcaZ8lvm42vgn3yNB5GNFB9LVX5ch+dBLsjmdQuQsye8D1ZR4
30ne2uxYjY1qBb94ZJQr1KW8hNXW12Co4DE5rGd7tnrzOmKAAc9o5l3Hzzn2jP9kXO/izwcTlQ28
UygpnExYOY/+RihUHkErQ1OOqIMzLxa7lMq4ZlWR1Ji4zhlkcNb/LqVQ83N3QAwMot1h1tUZaf+9
bA1bHzcjlB+NKso/aAlMG2BPFLIlncU0oCFUgbsdZ/zxCJLBhzZWIhE/F4JR8fYhTMkJT4MiRtJs
o9R2QttjIgZwiXVpd8w4ivU9g1RgV8XyL5m/i/WKgy7lPN8wXAWe3+09mjpJ8GivO2CpRGKwpm38
Q+drxgJkzO66CZrb+D0IrmZErERW8yAVfyX45aX1FzH7S/ATi66KlFLcJ7BXbPY4i9NW9e7DDCaP
h0uMqNOTCN3kAv+ajiSduo2sp7Nvsv978rJYSxoHtnZzpnd4y2XrPr2zdqPQ1b4OLXBYK/ORhXFZ
KVRSnmUMag1XyXqVrc0RV9ask+f0R1wp0bCRv9Mq17Kr3ptDiVFRieLmO3IHBeVBsHAHejQIUa5M
36GcLvf9KZPdB1fsrTZpyBINcj3X9xUHcU+VteCJtvN7wL1NgpgpTrNFxAqM8w96ZBVS3aeAxDSf
yw0AdMTq03T6VvzS1yFQnNXuFYGY94xDZ6cTO5EmRJVbKC/Lvl5djTPCaWu74jvBJnv7d2zsZnlA
BvFGPStMlhjHHuiOhJRMOHJX/tpZ3LCbyAbod/Q0rwhVcB3gSg0sLEOpXEQjGeiphFn6p5tB4KSs
QSI+n0NOJmBX2sfIeYiFhzy6O40Fua/PnydbojTgIupihBabbzew+4o18dAH/fScc0uC7M35Chh+
gld1mX25uMkC4BpeVcEzF0ePuVGyf6Lx+gkSeVD00C4qyzCc5NBgDNy+sHcqNgWG5BdjGU/iSK9m
9ceTft3HqPWcMV/07xvrCAsHg8QcJKrX3KtUASJTzHVdGEIlKsNNrWHSXj/rLM4bwMcfjZSF8utm
/aSxLDVhhY7IflUBsYiVzs8pRKVIoBFvzt8ZK1TvNWmKHpwQ+PFckE9mk2lLP/uAStdkfhvnkV8X
uMfIKjfbuzWq9blEPJjrIf+OOoqWMWRSQqgv3JE2KGeMMSZhGT4pqhBUYbjtjldho78AeXyCJIGF
IV1IOWnLjm139kkxC2WcpNil28p/UQWi3PDVsC+vwkHbG8iQXpizK43AyIdKJyWZsDSfI0c96kt0
NnoKF5e/YZYcTsP9arRu6h2NQothqNLiVHHB2rm4narohm2ArVjXxvKMFqswxDsxOttvWa77BvgP
sss9hOcutYcTn4RjYqyx8+42MI3OuYe7emGOyREWn63ZhKoWhcAUy5wPu443Ma+qycSxfXPHYwEU
A/1OOaYUAV6UUiv2D9C4yjG8T+BJhRW0AlWGHuX3KdyxsaAeJmus+e3YqIY2VrJjMSA1jWY7g3xa
mMRYqqxIv2zt43VQ+bkR7jbrpRHtvcWJVXgXkMwPcX24fGoSnKs796A2uCV+xk0lLVuAl8bSM/3x
7hFHcjuE8+lqmZIvy4rqAyGr7QhgIE9+goSXEbIGsb5MNzpV+qu8GG/h3KUZGyhtHeo6DYeX96Ia
IXbqw9YWwWLnUQa5ZUeX5SaYTwph9hiuk0nKAzobBVIFwWZdkKU2w/K+wSASB94oVleG3RfkuFrb
akU4pZRUdFeHeVHow//ZFylNrzCZQpzRXy1J6lC9zZJAIchaudCBIrdymAI0lrGH6S3F79W1wr9e
x4+F9W5aAXlHUk1Ka2zKvL0X0vLRbdZLTMzTbuBB7lme2/FnAEpoAiGAJCC0lnj7VXUJyzb8fmig
/bNfo3Ep7H9yUfymHwmlMC3fYhZ8+ORflMIZhnUp9H0ljG9VFAFd8KVO671U8SPdGoXQM+RuQfkx
eEZatXXF3jR5I0Pl7QlPlLbYLJNe8BPOW55d4fBLIi3hbQPDK9C82em4UVUKiKFWQ8lHKQGGWdmP
xCAOnGzPClZR5RcjS+z1Z11FuYDVwWmFY3SEsyQEQgC2A8YLIcDoKuHVbbI/c/WYQh+fO86KS+tE
uWuP6CDJtSQHUGAton0obThQgH1w2EccKbQCPkxI52q2U5zqpaEek47CJXP+k82frZ1DfWjb337g
hvI+I6noRpnL7VrLHL9zeI5h0GLN7VyI/jv7Yb5mbjTJy7G8rBjj+b16LdUoTtDydj/cNm/6NfBp
bxbbTeIRmmpDh3RULLuVZTZh0hBipM0uMV7x9maXzBE4QYGX7CDSaVNsTbtDYLH/yFYuX3NJ1KbI
lGSMgIT7NbQe/3iVfzDiP99JuX/vjiBMPTAUDhAXgxOfVlVB8Ufbmy4n+fCYivwdwSfsfMnNioTr
oGin/FLExMMi+DCxp+VQbVC9EvgWrDxqxsn/C4gdhYHQPgvAs3HdaYyGjheQY8jJTARTDQf/X7V2
NHN+6BogcXobxvL/cnyWnvXF/HQNqpcW3n7GSczVW0iLTjYzLc+pOOa6tvwcrThFwGV6AORKGs9l
pSi/hXyfItQFjuGG5+D3XM+SIj2oDISSYfR+xdT9nqMwW8Y5YHncQjps+lUa4jPXn2p+lZqgZ7aS
gGmnDIlOAKO1I3upCcfQ3cpZuJVioV3oa6aTv+sy5NuK2D0ArY9HFzr2Sd34Ab57v8Pp9VuOdPGA
eeCFVLPTq4ww0+9qYFgJHwiFOJE8ba/wKTDTolQABI5a0rFsCKRV76DpyEF1VsL50w/cVQ9w9GtB
Bez3xC9MfyWxMRIxo1ueKaqgf161htW5eeWrmVM3wBOPm6uNpIr6yXmoGIDYE3yKOssfycWgV9gk
eN6lbEplWdGRO4T1SRf/p0ckjfmGfhz8sdnvVHpJriE/4HosQCojfy9GlVgQzPueEhd/fdIk5h1R
+6TYolaRmRPDpU0UB0fR449hHSmuaHt/2kLtFknN5KprIPPi5Ig3GjVW0dHfahm2dUSgiUj8Qrdd
O22tZatBo1FwZa/9jKHig5V/jZlYE9VLQu8DVIeYrdWn5SeMlXlbQ5LtgEDK3X9UL6C5Of5P7LXJ
4eBgpyuc9QMEJs+Qana/lHujHS/rSXsQI96qiPHQGHNG3AL7UvSHgMxuz3ODfB0vW5tKvdpLD+9A
eAllWqG6haFFw0kX6/aQ+7j9eTryyh6aOQjubvPDAPkLgl1vMM6F28TBjtK+9uBWKZ6X6bFmnJBw
GLokjt1hNJHLh5u1j0rPpZgV1NI95v5GpoxjjKgqdXELtgSLLMQ4+pZyt6Lspk9Sw5/RtG0+TQF9
GEmbe1yrIhDlMjI2cYCwStL/5ApLOCc/oMHrZYolfCNiF05gDtB3liAAzYJCsDSfKOFEl6n/ZVHa
SsirTifMpS2v0S1ynMq+pBk8AEh662GzvNtTUNZaFgtMHdF9Gtbz9sFeqJQRaM+uL1dyvS9JoVUI
/M3sCLcjJrL7plcOBEHPTfTbWtwp/D06nfjP8HBvwMnCZJo42d1OAeHOM9YS21RqTUoeV08EWcsx
FSkNF0RIoFNhXocvtMGn37IzDYDPPOqECqr/f4mjw67sgICKg9DlKbjEN+UL7PEWXUA0FSGCkNic
iuyFnm42AWrh8Im8ha08C6Nyw4suQLBoP1+x/9wN41abKqyMk4Kg6fcoGMhsalPbnm5sUdlmKxqd
DTxXgwK4eIOMypoCqcqxPwuU+06MtLMnt1Q21BS0+aOsIF0qP7rrrCmu4yhzabuKtkcb3Tcitxyz
ISsrN4V/rndGkzI0zYqXDYYLMXvPjEy3AV2m38+Ngm7cIr9UfBeAb2gM2/LrgvOj/Z81STWlt+Bo
Wf4USTUbxEtQwEwAm5fFvqv0yUz3ZEStNeNEkX9nN+taoH/wXE5PII6BigApnp66TvBaxKOTLb2G
2xFQ3U3kB3OLJ0PbQALFwJQ+NtcO0wcdSmHkDRD7azZmqbff7N9Rh7jbZUoD0VzK504BfJG3Hhy0
2VTO4H6JgeCa2Jbl4FECbjnB5hsDwiKOfZWZQGiw7uHQ72Y3C3R8l8cAuDEpaKjyudQE7gTcg6As
rAs6tdZj90vxqXQ8TptRC9S3P9fEzcy4Bh03wFAeB33rF7+3lW4uTAmOS+HT92urQNk/AihIkvt+
yhyB0qHocsGuDWE9q/GMLUfaG4kqJjYlA8PA9soSpFnoDddOfpoREpgYSKwli12KeMfGFIU1l28v
7PfAYzeb5J6IID0PMa5q7xPWpeUeSNyIumtW1MqTbXtARdtONwCrGjP9NZdTGrctzmxn4dtGOBgC
bKkypAHUS+c0nQCSdiJz6zshp/I3PL/IXaonV/1y/J5WlhULGfpy48n6uPSMJ8gg94nRei+IJVig
NzRfOfFBaH2HFsEHmtYsITtB237XnTpmQrfX3pqQdfhOs8hLDFfmOPIaOzC8e6VgnY+q0PjxAUro
ap1ZetEtGLIlTl8iGaNTI0xuyi1oREfmZ7qvnonweDfTsR0X8pzEnA4kwIN/7Juv6HC6uEQpe/c+
rH4dKuBENfY212B+2z+gAGIuVGKGFCKNH5NVSfIZUDrjxrMn3QMjBzWR5Xmabuw8f8cjfyC6Vtli
ab/S8/5zmRA4M39TtJKh2AXEJevsRTwklliw6PEUibZ8FLmT6kIuHB0JMEDrVNg2IgQQyDbGCqjj
hXc0hRN0+kz2RYG0BA7YKl/tYE6gOBARTCz48/hCVrn3L3pue55MQ8ai6YtRMX08xKqOqtHAm3hd
4oA0Af+R7H33Hs0WDugR7OcLxETmYVCyiJICNEt22zztqvg0R+JXAsMaFYfCWzLO0XTfhvKk4Sej
AZ1kMzwCPvSjD9Orcfq4vX4sCtuNyrkWgjbT0nR3kACP6qjYuRukqU8ZSfDCtPIuJviSj7OS3nK/
lIaJNIJIQe1JVzgu5zPGpDER2JnI4KoZgeh7WaYlRNdyVzCZgxpztQcnwZ0FGHVkKCL5gv8AejRD
nkm9v/2JVQ0KtJ/Ufb6/NRK3uQVXm4JFy1846o/liB/GXZWkZyIPDaXJjjgY1Px7NvYGrScP5jhx
ZCbzvd3l5Tzl+Bx0xK7RhaGfv94xv1Co6yvJh2ATyGfiJSMIwGzoEk/WtZn164PT1dNaHLo3AkJF
ejW7XBK2jgSvUWJQJnEp6AAT92LKsFy9COZU5WvDpDbM7gLopaToB3FG12TDnlrUrdhNeicB06yU
Pv//IC8zMUQJC9o3mQAHJLooKYwXXFOqJzO1/YENumRvJfkInwXG5bOkOOtfqC6kN0Idv871oUAR
bzDhGtOAAmFrhgUrnToLTDnmyv96TV6HD2CwrxUl7ObgpUpsAj3KiNTmrHgH4j+guHnMGNHdDgl5
qPU1h3bnGSvURB4InvnqZK8zRIjpJwAUfHjcTgVFgRsZmzU6lkYewN2V0+WrEjSU7936HrJjcwkz
gUTqyP7l8gEDWG70IWwwAOQRtT0hZZgL/Xor1s8Jif5xH8RM2YX7QdeS7C8gdb7Z/Bngt//tZSqB
jX18RTI/iAoqnanTFldXbVv/mg1fisP/avybEsocFgDsuYYzvCAxf/oppuibPkJAEqfwO/1CwmuG
AG7p/PyD/n6EIaOI9VW5Ttbdn7F/Ztuobn2O6SS1q7our4OiixkNzGIX2taCameq/i4VAoLFDt2h
HU4XvUO/WcrS/04iyfN+aY6Giqglc4b/19EoDUFsEB3mU/WTHrL6psPg0u7+e8NLiJ5UfUiX18TC
ye5mLR6lLEe4kBkourjhe/ERyReSdJBIh1Bs2RjStPfWZkqsIfVBpphzRcipg7TkYKdXb8PdoB5l
qL11JGwY7QVPvuFGGlk9cP9g+APgP3IDzF0Fq4+L+a6f6vIWpBkuJ0Rk72uCdTQTbU7uA1f8/GJt
K89t/cSWRbkpOxhqKxhx437Oj+NqcwXoePotgI97CJDao8lQChx2bOrfkrYENqCgy6Kw6Ju7v/wG
JWLyXDIG8ZW+sGum9nRWOjlHpTjG3/x8z1u8d/nImEj6mWZ1tTZszXAG5lmSopi6AazR5DAfxDmg
u4agXTGHzj59bnS1zEvlIJGogvh2AsIQeaVR+8be6il2uM2d1WjlyopxyRHdRkv3K2U7AH2pUQ4d
K1xmmv44xEz0avJ0moCrhkO3aGmKlRKXAGizeHjaCdCqN4VtJbfy46gfOhV0X1afUlajNH3qfnGh
32HeYpTMJphtcn7QtsWVosMukyXd734vwPsDvrgdDt2dk7MPpKEb2Z9FpdroQcVosHTwmNU7dXz7
Q/mzGHE/P5A5V9ImXbGZ/4JdtAO0skelYXcD+m2/FCzCzmVFzfU18mSVand7PuDbz4p2THwcZf9v
I2Re48obhOQ5zQy67BgZsIBCKuAKr2+vGLZI7alAluUS9kZqV/xV4HzGXvV6R0aNanM6xRcCSThB
9LrDOuw3JrJ2DFzxBc++Y+AZ/a+QAYga9MMXjnObPYdlIHdt9Ot2DG4523/a4i0gZ9vECQuJJQ6F
fpN869YbZcWmZUtkxJ3S0KAy+96hP1lFGMF0uP3C93M3KgFO0xUzRFPR9NMVnZJk2oWdCoMFmvHa
1Dc82hUvCkDWkv+x9EAz+PIVzGDcKOBblTplLxmd+S3e5PPYgDhT+n3QPwRv3OaqYxC9Ve26oObL
lGV4sz0v+oN1Qf5XpU31vmYlh5jfBGF873Q4nvDae9grf8HlYbAgzYYVBlRDAZrFLZUW/OtCrovA
OAscCFNDgAJDxlCyClP6jkWTtS/Bc37IlCn5t6d/opFmThjnkGCjddytZu9Lv8FTeq7suFKfEbQv
ZZdXw+8OnIJZo7ejGtQnvvrU8kpTM6ujDZ9UbMTQclZMlanfK8ydQZ0LTbh7bod3gO5EZcxdEjk6
hUCATBjzqPpVz44F99TgJ8B8XyUsyeqe5Onumd2Nc4FoCjhJsYrnSf3gEhQVag/wiAdHPSiS9SCi
XEM8a3WhpgLJ5s/3n+u0Yx7XKy9wbViAhsAPB+MAtn18gCPKVoxVtqtYn7Iyi3KN/joEHnXtEH2N
bIuQkevmpDNRARRoqJTbUrVdBqoO1/hA2nhMEk9nfzJAavwn24xM8ljH7xmZnzCWIsAsMhDUOeoI
trW91PmQTJIoWKU9hFfKZArhzDC0elem84MG58r42jE86B7BBPgrZyJY9nzB++EW4pzk7KD17YRZ
PjSSJRCz+qu7tGKFLTzfLVi5D0yt7TnWSvLf1GEVbt7T3Ve6/oz37xpxAgj3eZ4zi3MFCetk79au
Nbt8jdDD7aiVXK7A8k0odE2Gr0uaZCAG1GammUJxRe02fkCh7wH4C8OTv1igYwkwhul/YsI6MrHQ
++oOm3WoKARyNddOiw7QjGbeKHo2SgLkW/W+B8ii3W+P0WDrrr1Jc4DmxZiTTgL6GwUjdrh+HWML
tV+6nbid2GHH7XC9G5nDh1HGroTxi8wv7KG9b6e081VJQbbGkqDlacW4/v0y9XjqP3/gylbKo7jB
P3SrZyP9TDX1NRMbDyYuzTTtRBrnuSIbVPMydyqLW+xW7uVfR1AJMtvHN8sor9Bq5GVxw9qdLZLN
ySC3h7Nxh4cYbZ3uS6AweoAxjX/uEiY5TfGzOASSVRD3jZpU+nL6G2Hqp0+daYz3qTG9Jztssh6E
MYyV3KyzEB52caf2PdofUqOqAbSR8CIcfK/c+YCJrAYNLnJLgq4SFbWLhwbNlIz1u/T/bJj/7ury
uhnROv8VjRgO5FDSXfrBZatCOs6LVQaXscRnauNsPbiVGjrmk7fkUByeYOZkoinpdfCO/5KOU7lS
mQdJuRP6hBtzRdFyfqoP/NVaV6gYuxai34fIvANVZbukaLlmbK13fYj71te7z9+no9QnbVHV9ZOi
SseOlzkwlHEPuLD4q5d99rdWbbTLJomlpknPeTN1Za0hL5qJKJU+5C/jQEDl+B0wYyITuM73Glzn
XWjeAfoW061HwXg4gPhkm6vRWpF0645dxiQbJ9zMr3aVB6aTVzHDMGH50byYN+pCz1A4ydKRp/LC
yEy/AdN2SHzjGOEl9lAb9t80pti/80aPfzFlwOM+jgnkZRG6+wswyuGYskwdjGZJdGRafi/Fi86i
EixSJFvVMsqmHhsknByO0kdfYmZaDY6pJrB/FwASZam8QcAzwF6WE9mtOtNKct2L60q8TK0QuJK3
m7Lfw0ommyPqF4jGcalCo4I7hvsTLqfZCLPxsbW4dyfR8u8IamGH10e0Si1ISR+2lQ8tGBUY8ZTx
enZ1mBxg7Y9PoVuGYHVfHuuTQ40iZNkr6kH7mSJUgKeYlhxLMs83jW+5CtHEE+QhibinYkfJkB2G
Iz8QYxpJhqgsKwt41kApTux4w0pak2lugG1Sj4A7TrjbSrSotqS4Ier8r/6XhaqjZS/0Cp2e9xB2
+LTTEi19uAZdLoe6KmpfDnQrL2Jox+6njWIYvo+gmGcWzeYNFUGFOAqLIkBS5M3dIBhrTEIlZgZQ
0LG5dnrjJpMUrnxF0Xy120uelBVV/MA3lwO0ur5kzderJsbLhUVd0yPEok8OBiy8DkNySKKEEqWC
erCPYcupigfqZo0hHWpK4OCGkd9PF7IulGtHpl/PSKXve4LS3B3P6HUCgH62PNeoiLNFnUawP/dJ
KX60BPyu8ZFtfsgm+51tEjRHu5CKlgBppLdJCEXc41eJrMn85RrWNPQ3ZzdpMy4Zi3pXOMzAv3kc
TaFvszefSMs6BELqHMPGOJ8b/ikktZCXw8nb9K8jmQi/EPKkEzzEx1KPG093/JkGpKxVSM2yL9ds
hn+iTJ+8sJNt5pNRtX2cVTM4IAvaYgneZmaGl2fVRzNt7JIMTet622NEguaPtsBz+/Ce/xkMB/lY
OWMOLnmjG2b9s6MNAztEruvGsqTGIWE+FHnRvsyKbqeAZLPTQH+CRYyPkL3rw4Rd7qA4ePmsdWLk
3J7oZJ9DZrxf/Z0fffkcNCo2p3rR8zHPzH4EidpkU9ngAghwi8k8RDN00UG43lHZsTnlxb+Mpyh1
5FU1EB3CW4cghSkOacd5Hwp3ZWrx8a0jPdaVq5DK6ytgT5J0JL49CxDyUy3vykK/htJ8TDgsMdhn
/eVIDQ0ZdS8sTDupApA8nyEAbB9xlz0o0OLQM1MECvV5WO+5WRSVenfv1xz6OMPjL2MA4SJVR+Em
Gt5a4wgzHjhNlG27+3wqSRNEXKjXYWsKcZKMxi3Oo08DjEO5/6PHELh4Bmyo3ug1XGBCuh2mY9du
tGH9qTtjG3tL9WtLsOgMSHJHhsmXUUwyvORZ5xQOyi6FnxAKswQKF/Yci/hWoE5jRRyvQQ7Nhy0H
AJJSMaeUO92oHPUbROpEnqrouftXHOCkM9JQHCzDuESiJGe2KhjO41UerD64mA45LM4EGYqyhaej
/85Cqq/g1558CyFHaorcx2TgrwqfwrcmaBNUYsugbjVUseJHrPed/Es1dhF2G5MzTLv86HOLRNHG
It72wcbyOO/GEb5VAb+/fL8IWRIEKVSya03rKxr9HaTDDLy94G3672AmaBSq3Pt3i5zHggcnmA2F
6nerOrrqwDtW3erOFVmGT9SzAsAXeSMxr+1cgIpKItnMNYUq+VoqH+Mk8aTPHalNcmygLaVcJN2K
yXSUFlWAeqKb2oAEoDiy52T3YWFrHLIvxGi2jZoL67teOR7CHWkQqfpe4DZAMgMV4S5V6CJSAdWw
MxlFq21sQitVNbq5zJ/F8YqVCqXPvKTIYlUdqvn53DGAdej28FP6jyVpX9FXIwEUmLiATWeqQgB+
yZcc7V1v/lVCz1NSVGOpBKsf0YEpL4XM/BOIFmOfbm/Z1mO6FHg6dyjBsXxYDmHgFSchRO04lGLb
V1OIHy71ohjoSJWOnGLwD6UxK8OQvaxXPb2KhlZQAXGtdVrajtBPLiAoJEW5rRXjhIPvDv+ZHCy4
2Nuq/H3LvEGCi3kAQIii07cV103Mywj+MOgRYjYfnaCClasI6mIcRheQjMpZkQSHI0xfBGRYvAjL
LB8uU0gDtPN4Try6T3KS4dIbcQuarl3zBPj1u30fwzBjEnuu0+m6lfdgJJ3CI6JTyZH38ckGmtdJ
zcISiMgIIui5W5MOuzXoBAaPZJjdLktMG3sqMHXBFQdRfe80SZkFXmHD2y9Rc+eynjm8XSwS6hqs
C40ok9zBsfS93vNR4+Xp8eGJ3zEcPO1e12W3pGockpDkENNufzWlR07cZvAL+RqfOTzXBxPoq+/S
MabFNlctDpJeeuaI6lXGQsgAoV3Zar4Jgp0Xc7I520vYA7V+t8/dLhsUM1TxGik/FOdiFP2vV6yA
QOJO8ckx+glVqjl2MOUY6FvTR9owE1WW2vFq0QZlX1jMHVKqNfJePLdnF8kHL/kz8zAKJAGh5SYJ
+G8mpSMae4Kr75LlVuMa8/wv3F8U3ZTIP1ZDtgj8IEJmxu47irWITpq8vvL0yjhKMKNKeVVzu7yV
G8DsGkQ35xJYiG/5FMwPd8gBAhOo8Y50CPmVbTfqkxAMBoap8HGWAvHmRQMBEp/ZsqdgCnuonc8O
JNinjY6L8iPu4TzCwPcJHoQX79fCYtfkBXmdbf5HFeFPuomNLzfFdpMiLoumMWslNyQcNl90Bz04
wK6UggDKABMe5dWmbAhCH5dulwzG7/soJI6sFmIghwW02QkpcoQRLs4usQjQWNwdLG4hyFCms8HT
f7UjIVfgnux22LgMHN8SzCXfZ2Z4PNaorsIRZmI3FW0RVGRH+A+LYpK4IbWhLdxcVomj3gheSGKh
hHYjrhQlstXniEWZnhGk9t+FbJGpxHcmOg48PNssXDYSosewFuuIlDdFLyLoNmFyESx9/DrIImnb
5ujWPGdNDoYvCsbt3ruwu1/rF6NSmmfLhOSRyZuP+MGJW+BBbWoMTedV4KpJ48NmuL2PTkTO5lUs
lbDGBImcEMZEVRBBeLHpBVgj8uhD7AwzKLQZWdQ7jgUIJcs4coFhT8sR5SdsvfjmJn3jJOcPenaT
Ne9wwpY5GFMcrbLExMBaKxRVvMxsF7GyrAKlVuuwwtlKxfm8pyp1DAxJEeDF/dmtB0LxZ06UK3qz
BmEMgMoKBLH6XF3owHgSzEP3B/E3J58GxxkO1iEfs7ir0h8W7QUG0pfknZ/O3pbLwaID1Ex9KApZ
RPCdEDW8hSWS/PD5RdW1Iwv1WgI5cuhG2k47vLnlhwDbhpIfFQlasRlGVCorJQKh6Dup57Q2fBXg
JK9eBMoEL6HQaobjC8GnFHpLK/YxF6A2709em0F9p7voi4In7ambhhSUYKwYVo5lvvwWQpZKfKbm
Ary4VHOFFFbqs7S1nLUVtK9LSpR3SznB7srIPgX8SnxjAhX/dKUP8gRPBi8cNIUme1mnQ1RcbyP7
mR+DNltz3sS08HZFy+EOLQDReFPFA64OZw49ifopbmwO/8s9jMt/5R3uKFj8H4Cqumlpn8M4GxEt
pRJF3rklj560txmM6RXcA3tjOoUDI1XZNxDyEQP3Al2vu/rnmqr6Wn78JQA7Wcks4wWCwRtEfjYe
uEmkfMV+iIiGwYy0Qu26UUQhRZfPVNka+rW1Xb5pTf0mlz/62QVrEmAIk/DEXqDnVWyM2f3bTM1q
7Ev3obFuO9/HPZLiOlTGPJ2RXWq63I/oId1Avr5I8DjY2iY7rIDALg03gm0+mOywyesSFpjPimvL
xauvm7oofLbgJSH6E3swPtbD0go1EOLFCqg8YYZlPobql7LNRvKZ6/Cj0TfE3YQG387p3SL1QJfE
4cMATv1WShHbyDCTXMBYJuKTecSPIzXsItocVga64ix1U01RH9P+IOx/KeUrJvxEWO8SRyKlqkUN
sjxoGNw7rBfPari8a705UYDXQZJwvPcemyzG6X3F25qtWVe7pa7AtLgIhFnOx2HAkLLFsWQfXCKZ
UWSisg106FgeabpWHM9tnbkcPRyLi9P6UC2z2Tpr2Ex2KZiwtQEiSnqTreD57tWrOwPS1doaxmrD
pW0x6WXiDvBZVOjCbgsAmUxbiONmphF3tJg9NTANuqYavI22LBQqzlnCpp6EhOwNI7mRqSHn0vg9
Au0NkDZvWW4HRpk+glv5xGSazYL0vvpqvxwRubmDG6x64agL4EatJFr2i4ons3hUtPfxOFK/nC0K
iEdfs4C67yaoXr+1O+HOoeDuEncp82WdybYpPzvru0da81isKpO7cu3kLnY/u6XoGTXqDXs5swM7
gyPcAiCKcA+MsrGx6ZADFOINld/zP4OeVygeRKiV2kmIUA+wtlr7BmMys+vkDoZCxaCLEmvNad5L
BoR4782rrUTv00+6lYK2tZ8kJnPWOBaL4TuBRYgF+MA6t8NbEaX2x9Q6F/cV4V2sBYlh8wXBgTWx
pgxASD2hHi7zFwMLImslCznRrZLb3+wP+Hhn2FRSE+S6ivzmLXQ3cf3TM303BP+KPAMrsjGdVK9s
CkNivQyRyC6kePjkZa6JoHP/gu/0hbse7Nf4WDf3fC3mM0Ko22o4hTc8mTlNcOSi4s/LiYfAH5BF
uPBAIzD+Z8lFDu7WJm2AJDqp5dpc5DDpbHYyOo5PlSw6qMvh+Dyo4lUhXZKS1flSPkpUwLKK2vYa
8SwFNFMqd31x6zNzXE6ta2BGTjRKd6RvQI3Ln8MyU9tCz8e0JhCrKz10aPqdv8JCVtxKsUB5zLAn
yS4T3Gu7wgd2r5SsIEmoNAa0aYP+dUFRqfkmRSyMtju5MgLCUIlb9+AqtMUVR0MKp10vF89dw2h4
isaZCeK891XvOExjjWyKlXIzsOchBgRG2FJ1Ly2rMO+nNkTILH/1p528x9Ft+l04bWh0g9NsQPvm
zbeaZAffZKjOzGgtgdNjIaQ99HgoZf4zmFqwckiwjL2pqYeBVSG0eR7yk4R5+ri4LjvYoK3DKLgL
Gz0tgyO4rfcR2EkHkFW0U+6Cs50BQ6Bc/lZzdH4JAR1L1gpvR6HzG8kVWsP01bcqOZd7cuaMBVaC
nD1aIwznPqdoM8g49uQZluwGpFb77XuTOVGYVypTT/Zc2ZwRBaD8PWOs6GWLPrCAazcFmJyHt367
1v3cQjfL8lUw1dNIYr4o3Z7bpo1UpvY0KZY8Py4S0rMiOycVpwEHApHM4NWGkQruU6GlzSTq5QfB
kHdi0qNrwyfqZafGUKyna2Lx4YTNzlGtZdFPQK54sv3FMBi6KNhztRmuqAsvjs2eI/Td/Y+kAJdw
3i+ThBsW00lu+9vJz4EiRSVyViAZ785b4ZaIOLPAyJZ2sZUCbGN6QNpMmEe2YdTTBgmPGZnC0Ivg
QnfnpSD/+s3eqT7GdSVBx8fTG/atmAOg/p+EtB6fFKb+9lU5C8QKfPb6iNkD4rs71/hlpVHDTJLS
5Fpbi25Lg6HRkujEsEH7CJ0IPJi2yiEJ/Yo0flcNSaGeYtvF4cAsAeJ9t+gCwL2q08Fw87sh8Pgq
Nv8Z1SXFui4vrqHLl/D4SaqQFl0aYQERpR9k8uSxVs7n4DhB/l88WS1opGeMmkkhwh90WN5zd4f2
EqpKJCc6UWwuxzyd2IwmZQ8bDjFZ09EqZzueR11l+JJbc0PrTTDTisQgXOsiMaIlOajk5+dKJxAW
1lPX6hTfGxouX4/sQ4DyqDvJnQjsiX5Ks5kb2Pf7ZqybSKa5bMEIrSVs6fA00VpGRczcyRGkrtoz
e0vT2C5JBktqfUBtIQdHUeLh3TK4bs6wCXT9Hxfg928EwbEPg1cH1nwtHol7+420LQrd7s0Ma1c+
uv5YftioBefi8QPsENueFmZZLU+VU+brUsUR+DCy/aPkSgVjyrrm53yKAg4qM0glWruWbdkJrlw2
knriRenxz0k32I5ihgqoypZMAyvLOIg8mXisH/ck3S052xdHr0W0QAL0ygqRSjnA1O/cJTsThdGn
xSlrktyIp2xNj6p4+ocyy7OS12I3qAHHo7yrPkRipNs+9iwWyWX4U9l+JJzFE0L/iGdtWs6n8Mgu
eVJ6hoM5j3XABJYfFpGGeM7CtFNUVXvgv9ju1YGIe2mVSgCEpV+iqCG38j6xTU/3v6ij3WfkOVZs
8N4n0cD+JiwoJpTCQZYLsWQiEtJUQ0b8RQb1x/P1ZS05O3kqCXvSkSMen05TAFv7qCV24jzzv4L1
SAAwEOsaO24ZZ16AGoFUt7yGmL9oQdYBOp6UDpSxiau8HT6X00GTzGpEPiRh7nXxLeavIJITeB66
S8dfidOvkEvwb+E3JCsEVwDpWiFm5L5ta1SBKd5snIHTF5Puk6Xl4uWvoVuvIl+Kq9w9eHjZ+QiQ
czqTrW9ckYjiBBLOuzqsyDn9grvU4hfcb0RV20BI46eEZJDg9FNSnxxvBMdA082fiL+nRhAMSGPL
H0ory9ysrjw71Tvkmt22tTZGQTJd1yCP/7xnj3DNO6DmfqO8yZcQrILkUDHXZjYQK+RSbby2VPOG
xSXX1ik/KgWXp/mWe5LwQlYrA7MBa34rB5X+pJWFFaBkPsO0tuSRrdagrMj6yejuxfZLWID0blO5
uxdt8+DTV7kNfQ2I1qeszFXIE5e1VZqh/jFdHTsM+YVTlEPZ19qOO22Usgvf42ET7kykIGdPfEKp
z3vceGzL0P+Yj1EgPGbJJBDiCjkfkZkfOgBnx6KHLz+VaLRc6Dxr9Xzrib8mTK6A7jDT/uihQrRw
RRgooQyq0uKR8OZT4ZIH08k/ciT0uHkKBVXaHWJNj1n2qwc3RZXutOetShN5CWQcPvyFrpjKBZuX
SPD4tm4Up9ZCfrXR17RzSba3yGo9i+KzQvVaPP/NeNVuVwhqN1KvTj2HdS9PuxF4MyBr3c6qkJ/r
Lthk8Pw8YSPkD7jI8OGkDKBAJZGKf9HeLl47b448GNvulHiVEAqOhTua5zd/qApoL+81EAfXoOF/
mQP3ITeAu12fvf8iMjnpUwqCihCb2o7M+bVR+dxAhdIBbYxw4QKz9GxWSDnILWuhNS1sSuWrRu5Y
lpUTaoldXKcsiedDYJCsLk2BdJmr6jE0sTyuhZ34kVw+M8qrYVkkjuFw6e/jPT6WY/aAilUAuGco
CTVVIfy1wCU36R7L4u9rIjU3/cfFcUKNUsryQ4R3wC9KgdwpVmsJIH7PDVNFzOVnnmzbP5ZA5pDq
y4azgWXb1EDho3b/Cr4E+hrckUNT+8AQbMyghm8katkIL8ozGNGyRrEdSNCd5nxxlxF00RhMjBy2
n+ndVLubzM5qRvn7Hxua10ffF9cojuqbAzlZaTaTVddKs+KBggPCHFD70Yw2Qi5d6SmDJDiWcVTl
rjjnsTktmPkirAx2WlPbtDbEQRmd5dhoJmhk2Sbz1T3Nhb1XXGzSDnWC/hUt502+lXLQlCvipxNT
9Qcbm1Hd9w4p7nLUEL5Ltbwm002OGuc6yKymbu6S+e7N5utCaGa5cKYA1Ra6JXktfjfZpMDqP4Xb
9rAMfSP0vFalx8eWZAmOTErmgQnFqFvru0/GgBtfjOirDDfx+cLYkBALrpeSe6PQFzu4YI68G1FQ
47MTnr3MCo1Uj0cgi5OM9lqLRoTlsyWKmNszLDV2xtFmkYdza/PNKbqNxZz++/fjmuKRad7BdClb
GPh3DfAB6SC3ry/v12/YmbVCCDWa21qKkUsWkx2/w6InPwKluMd+Flp0nn6ICqOCtYL4lsT/rkoz
GAcbtPPLYpYtM2vzWXjN/fGaTWM+xHXRE1TIKdHLNmSXvyIohigUaA5TLsONZIIvKBN/rt+aWyAc
DroY8fisu8y2uL0rG8hWBC/1vHPCccNyE7bima9TrY2b96nIz4GwoPRhGhZXlWYWSGG6SUEhRIiR
rmTYXZI4f5rM6aq7IVAzahwPBeAWXM6t0I3g6Ppytnkf0peWbL0seuDVRQp7m29S1ndJAh4Dzbci
spnxowXfC1X7RKzJwImmrpyRfeMZl8CbAibqXf+4SPA2dYnuMfYZRl/2zD0Mvuij1Vcs9P8QMXC2
IcsM9ilyqjZMYYE1TJb/E7vPifsIx7ppuFqn/oaKog1QaNqqqDk2/Q50HUeJs35IBTyIuVQD9XET
9jJmi1anLf/GrxfSZc4Yq5tlRohIDiq0o9WqTWJ+pnjMPrwQuDs0vjeXQBk1fpZ87BQ7/eF2gCTf
bIntD5tfkCkYgom0moyUVHck3oK7Aibu1+elhPjBSsIwi63BF9yZyM8VH6nKqz41xj4tj4DytYSx
CCNADo7aiL2+AovFA7x65KH/4GDYIZg0FU4pnFEeQQPRK2uD4ySqnleaca+ZasuA0N4t67QDrYmB
nqJivhPBrI4VRWIlCWJAuUVig/RzPgnjWyDSn84/8lIjPFcMF4gsIE2mfwJFAqz8wvhsyhfPgu0p
8WCgBXtRjU+WVaaWa1whh71yPikJfbzES7Jiik4lmN8lmYsf5nW9vpayApaubenZmYHDj2OfKESZ
sbRIq2aF5dDspqxwaWKie/dNjo1+ljJ6Eef05QCfFWHnvPhdQrazHbaiBq1z/Tik1WGcz58XdZ+N
wgkn9SMUEMVzHCgwZ9vXqYWiTGIoOVdRRPSamsFuSBQ0Uwk4YONAijloCPNDhlGVbXiK8jo3zwTb
c4SABaiyNkMfteqV9vsYORPfGNrF7kt5mbh21OWMkbMXJtOLiDznjm9c3zA+zGUYYsCEKKCOjnue
FfvGuZNWYR57h2H5FEg+CTn1M09wHHthv1EbylmYTsAP/R8Dc4xp6os2Q438VBRv6wuSI0nkLjb3
zdTaoqZp3CnHzF58DCTJuJtRNzAHtzfvBlSUNa8nPEyetNHqndnNe2U4oziuxJb+cvHYuxWrlJBG
5PnlVgqENs7K8WsLYZamj+9RhP+pril4M3xmeEEeeMy9SNnr9gYMAVXjkW7grBVuDUroVO45rhzP
8QBuWgzTC5IgTv7HM3qM4h7RllewH3gqeZE24kEYFGakpM7drSl4twQ+SwUYsY4TIpWzIo1IGNaL
0XzW0e45/AWWQJmbRqAQeNPGa6DLm1lln4SPjqqlDEj73GfnuWj0wXYFBus4eOZkGyVXU1HjsrPu
SpdW5oi9dZUWxsW/48zxiRYziGXSAnzrWsaQS2JTLsJ2Jtsx4D9a3vkZIAu8XRw8m7ShT8uN8mkl
lLVtIYSY+Lz39bsryDNOBhZyJnWx+FqcqbintYstf6/L4Epw3Il0lTSd1Hj/5G4P+QUAZoECH+L+
PMklsCCsvWpPQTzh5VWGycoGfydCgiq1Ymf+ffBZ1sp7MD/MIArzPEbe2HBf9ppDPXBalHLxhBQZ
bJFWkhUTM7dNezzJQz7KGbEVXMlr7RCI/nGDyiRTHvArRMyatr/fgR1Hd55oyKPAX2clF+HnwHKG
q0cZrZmEv+vBevPlUuOzH6YixAr5PPwgC8Sf6mBgT2eXs8inxGq82xsn/hr9F1zTsJo4NpGMSpSm
7pomMn9XFYGCp/dXeV5+P7iXJuoqmsG2fcuUyY7z9zC7rm7zFslr4WfpuH5x9bO44aKlXIjcQXvo
qegF16Dspd/8bbK4GM+P+bRfUzW4u7NTDRoH93/q5PbsHUxkH1u76PnOCRV0qFiDZki3aIUdGC66
QD+rU07dICB1Y4UDxGUsTjU7ga3iyFgHJoqhbBWHBW2QXd+AZso0aaBEZ3oFQneNCm2bO7NQ5+g5
IDlpAoy9nyzOQCcAFVoV4Zik4b7Zk8S4qlePKfDnYCUeqXTyinwsMVz9eqPrIs4ErrDHEWD6ckAS
TFBQHipV8P2ay0VAuW8JSdRB+dItF9tUWUHB2ZIScxF+59QQTJ6OfYPP6MtPvG1Tw0NzvDtBQTwm
Cyyz/OdAUwzN/CF0dR/n/B4jAcM/ykxlTiDnXCf6FiW0qKuOa9/Xfk3Wt46LmkMtYGCijcHbKheO
rlpLNhC2o7yqn4sLsdIWr2K+0yl3WRmd5su0AJXynxeApPQQshrCoQiuHvPdOS4+cCf9dRKZ6k+d
6YRKvFgVmmi6BAuYBQV1bUIFIdfolU7yjp9NDwCCDPrOQh+8DvWDRWA8OeTsHo+rROujtJjJFihJ
vQb3m8i6VjXGzUco0DGN1VCC1HruoYuBm5FwwnISVH3mpbjSB+JDQrblJXKA+NA+jcQBHt4UFkJI
7hHyHs7pY3u30S/4WRdqIx3817GSvxgWHOtN643FZ21xeQWOC0XInH7+8N/KeYFKHDlWIXq8mmC7
Rm9s3FXmHX/KPo1tCgfLRPZU03eUDZNtByhuqklg668YXDfZgWGKzn7TKu+RVJBTeRbGH4shrvI5
ABUxRDUeAbf4oDa+IKlX8PjNh/bHWVyaVU9HxpaahEhEckAvwUkBW5U6kDSGp/Oi8EfBykQdv3Uz
wK7CGvVELKWVUR5ToTFqqpq96A7hhpmOHOwVhFgYpJlPaTuGHdeI56YVkaKUZ6OlPfDwWMYQITjP
iOE/QXJxKglfg6I54DHNu4+t2vYfFFSy0P9V0uWSfIZqmTz8i1X3KwRi748+8jrvEl4BHWe5EgJm
mPaRf2978Qlk1NwV/P0zuVJQ+zUxQ0b/PgiFb7Q+CvFgolkwxFvv2edTxypj8oKjJDBgDkgiSD6u
inX5KiK561HbWx7OcLXaoEZyk4eqTyyz0TUrm42Bl7tUJbbF4g/KaOZFdPYqNfyA5zLqaDXGWxsO
u2Gxoc3d849H57BiHAsb8vAeF8hvdxnARTLAbExEOOB8vmmYJxJz7dz9TGik20Hdt5eSOhLfJ899
vc4mFEdscasvhJedGtfQuNosH7yvg4be61XpINeHS5b7M1n14lnbAYuzL6HIiR4h7OXDDrNBDB1+
fzs2kxIhaCXW/YcxApG+SO56r2kJOsKsWZa5XwsO5XvKB8TVNI0KDo/E5IbekbPwmpG9JIFyh0bP
wYBpiEz1htg3qNPKzXnUOn1bL7SOGQrBQZk4ZFR2TmrPwMrLJN2QgQd/eRCtuz5LASzDWsomOYgb
8PYphaM4u4sPlp9jSxM6NKU0unycEujZbvHy/HAMVHiE4DOQtwL8MzuIAg9bS0B/yhnzj0Wk+/bQ
3fNBxTWFrcggk2ygtFCiE9Y4l9GrCgbNZBmEXPTZV6aWwyFIvn/ZuqGRMogWctEUhPXyIr3VnV2w
Nx4drHFKJAaVW9qIWfUNFsKT3mUxfKDgBJb8aTtYGJNgYEP5PvHIyHIhKwLG5IsDoxF4fD/ntczI
DlHPE5+iFZdq0UjhWuPCRRN5BoxBGAdNCS1IXzFy554DypGzeSx6cvNP5TLLoZIbSSwTb0gI90oe
Qq8+49M/DfGW08CZ08M+lwbL80uyyJpM0YqpwNBrGM/Oq6SGOmy8BVS2Mvn7DCgy6dUuFawmlqnZ
zkeBZO2Q3QQ5nrJKTjaBOoTZZYtIGgKHgZxipbv5y0IhvmOxJ2gnTGrItDh+OUshrCZfz6Cbvpbx
LB6fF/e2d8AiJWxt5I8Z2ptU+QuQ2qVJ3fGmLNNGn/ROM3BTlo8L6alhEhMjll48r4WAKMQ8RHo9
gjtsKi5tqlsmcajVNxrQnOX500fnkJg17fmZoBm4Mh4hsk1HV5zd/XxjoZnX4MRF6CC381AaEOnE
As45R7+/bFrmnsk3ByGYRU+S11GuUQYe3Lg0PWB0KpotrdtDNc59cz4H8jhTCzhoba4sDicWkpjY
cIPzx0Lxp5T40OyejoUNqs0HSF4cRNQTH4aA5HpxBDfmYgs2HwmoXa0ezZlPq9X4H+xT6danCZ94
26nR3YU4xAirk+KVfV2fygGDcXEGsBpLXjm9q8MTb3ddPr1sjJPkRbyy4+IpVeUZYmlsxK31y4NY
03qQB58JsddwXmnl7JrB3DR/OSsEMbRsNbOlXnOwoU4QE0a9xqK0i+1E9nc5ZZCsmo+adTvpaG+z
bixL6v4wrHgdm1FWnWdVyYWPl7vMD1svACsI8NjfTnKPH+QO8r7DOf4C/xfoC09QXs3xDsRYXxhW
8LngtZAQ9ZmSKtPVdiokL7HZXoYCvYs04Br12WPXurPRpb22ZK0h+J8eHE9a0T4Kyy0TXnugGlAB
oTiaf2hHRQosGLfiSLek0sO2w7b8FUlcpktArKC60OVfnGK/NlFRlD0SJaO/jPJ7bQbi1FGnrSiP
wyU2hNMcn0V51S8W06H5T/jVpBtsUsWh18ZWN0oM0zvXoM+WzxYNQqTTb45WySz+0Rs70C0YFxlf
iPZrMmAm5F7QEJdBx2edzKxa0OFXaXGUsb/7w5PNMIARI1N3CKTH57PwY3HDTpS8B8gnwTaThRSr
9n2AUSJGxl+DP7GuxwgKomquJQI+a1nSQz6yPxF5nwU9up8moOz0iF5VQo8ThpV9/l5haRNJetkt
mk+dbj3Bu8+wiv8jz+o7fmVHlUv6bVj6BkSDLsSjfsunxlmY0flfQr3oG5tbLbRsN9N416WZ6j6T
9Y2J20j183YKhWFdK/JJ6nN29vDURHVFOY2cj9eKroHnXdehuep9MqVO/3GZoQlN9j2qZ9EhLuKw
BFHjVwlGsELgYn8hUXTHQoZg80jZTmyaxUGZpoIz43ct0UO+QGd4wMKdK0nxAIg3K7S+OkPMBCyW
tyMaRv3crYP8XB8c8WxR8ZkPNLxNK7VTT30d1Gh5xGRSUKo5cP6VlM3yylHs5KNjSB+hSj2XbQIL
0kPT4S/4OQmUbKVgxiOHxda+NxvjZnt5/ndEU0t7DMTEwN14zYJOzw5oejBwYnhAEBRfaHJJQ9Zu
toqJWBbIxKSGH0Ok5PsJ8c9z68Dfdq6dwzYiKmXBnXPsup/XgAIWeKWs3P4ygIOe9eqyb+WbSX5w
GXH84UOxagdlM6RdUF8xzYa7BFHFbam7+JovWeHIgmJv+dArpzG2a94/3ew1PxwKNDidkhrSQV/d
TGSD0CEg0OOt2vOr64gigzZJAE07gqcLPZcBFSx5zCDKY+wZ+WJqsVqchJzLeUdCVRZsajF36aTy
cxBrGzTSnblj8KHago4slJhd157xnSUD+/5HBo8q4HnDOcCkOygEGko51UypnazKElBpMkF4wOPh
YcPL8sqYQZW7ywuTyjOV68u6jZtGSuMHlzHND7dRTaOA6C6PzNHFYCTaXnF+slgI+b+NG0wyOjz5
+6000bc0nyhjLanP8X+2P+d3yRiJe9Z674al0PJpRQY6QlcSYRm3maycBK8V17Zz4N0q03j6h4aK
RKOiaUAPULu4h1RxX2009YfNnV5hwve+Z9/2QFzUNlxL4IqQybKwdCj2GNn/4rPLvXal7f7uzzOw
vp7o5KSqe9k9/1L/1RZrIU50/2m/m0vH/x9MyILldFyYEElj3KfgoumokV9p+B8lV75zQvaGMREI
ioOJhS+VV0Sx9fmq/U2ZHVmNj/UWs5PBcQ1GgcUbA7O9JobI8XCr2q1Uh3QtFnTlvO3LdG9Y3MMa
dzBa9tHMPgdDKB3Kd0lmB9QVmO3fLCtx1VdxShUJSrzM1e/Qo2EyPKiZF0XNEjVFQJnJonO8yPJh
L2zi8/FrLN0AzGtIPb+sKvLatJ9/tiLXrn963gLErrj0tpw8+6kiTPCW+GTJj26ZijkIp8SxZIJh
NoI33HM/S+9Ird7YK/B+WsFiQiuUh5jra7LkkHBLkSiz5OAOMS2ygD+VJc7ghxcAnEez5hYzzBQf
VSHSx2PgrX/JI0iawamW0eRwmFYwmMmMo8DJgveZ4blzWMsvssP0M6M8+TNOEW4McsW/EwSzhw/c
BC6WRMtoNAiJtWBiO+gdQzPC2D9fS09qTORxTyibI3QGCxAsS+HsT5XSs01eZPQJxImtkRcBHqSe
iAprSef50fgFHsTml2GvfAPiaE2/x8TH9HgDd9kRgINb3hpBt9ZHYZzCVslxoY40kn+IPaSoHelv
ZQmJQ2kLTdgReiBm99FlDepr5Nf5ZoFg1+47uShJgK81PXKy3NH7HRot/2Z3iwizjwX2dtwkTIUa
6A/2gBJoZWRRCpICupefXo0RrdYyRvfKReTWvYNU5SCSX873ZYhDeHFT924F5tOmiCZBYQGYX4s/
wD0I911mFPZOEg0vQ7lJVd1iNZr5Rwnk2vo0RYsm/LzQ45XsO5Qg/+yBNgmgLT+j3MNr8bE5584h
TVOONvOTkV1DtUsT6zg642zsvqkSIKMmTeWeZKVvAeYuhYegYxjl5F3vmCZG2tSOxdfpUlxaXq4/
sgtUqm/OyIbuVRWc2/oJ3A/nMrImDOV+eeCEgcSL9pzhT3jms302BEVHPc9fI1gqQZ3z7Jkf9r65
bS2w1kI09jDMkmsNZhx06Ke39Y4Vn+79Iob9f0oLID7AtwbeyHJF0Myu2QDO5fCndZwQdwNA+ZNB
kMAuIcwG4V6Yqk7IfPi9pvsDnUefTdMHLPf1U2X9UP+wWjlDM3bjPjvRfs8UpReyLckRyZ9kc0dR
sDyOlRf/Q3AqRvVzFwaFGn1pbhgupkftTvsFdJHconv0il6ztT6RRQyhoxwjuyZlc9dlNX0/cIDO
GMfMO1jl0zP4tNWimBg59Dk54LQqO/LgQ1dV7ezjOcluBEqK9DhxCepxJl5tvNKi0stqfNPY3DjN
3UpGztcs8QxfZwWM22JexZSxcObUbfNNWTUY40Aia6oHIw4gRLvmSMWPq38YNfZdnaVXSrPTEI/1
h+vyJd97IekczjV+aIRAT9/Af08uU4zbyUuEvgfgEbHvgkX2hfDTScQqtvsxBJZ2kT5NIk8CuHym
URVxQHxeRXhneKKlVfXo+hYEr/T6uy/ACOidGp9+UztiaFEvgxyZ7t06jP1I5bAvWVwwtlDfZK6P
p0T7hPxD83Gy6BKgYLUv6nuwwm45RvkJk9Ni0NEjzoqGDhdh5grvOPPAdhA1/J00mbXpJ0kUAlEy
WlAaJFGMscx2//J54UQnKx5a7gqderaA6UageZleJmvQjbA7PvHqnH4o2qn5ofjAtTAhBkY/w697
JwXoRQ7JAb0rwSoMg/3TN9GO+g0TSzk6uPrZfwDaHj/SKhTtFWGW2RBxX27/QHvuYL+c4PYKZbjX
j9vB95hIWW8fQNh5Uq817hA/cKt1M9PWqM+V0mOuQTrluchl3WQVHY78uO9lwMua2SvEjdgC6VVe
3fPD/1yTGRyyqdwe43FTKHw0dLil2WnSQiDV+OBVt3wgqFLUtWqhwA/wJtoQvRuNIF1zf0wszXJA
SAMNr4YNtPEDAgwazqzHTqiJQETik9YXRRg6Zn3DmG36BKrPcXzMHBQ3aO7Ghx3qmR+q6hyDbewp
RBDK3sv1abyJzMtK1oBZM/uOsKBkRbu8+VajGHjsB9E1Y7IJkqiv1/uhBE9ml9VGt0Gndry0dfWJ
qCwmJsR1OOENHE/2ETAs2HGkX0T90qIYBwvasvD/LXeneq9mKp5mJP5UniZvjtdqzu7ST5TAfTMt
+KbRiPQ7uNOP7JhF77/cnor9k4nTBC8RHU29FuM3C+aREuRC7/LI+jjVoX89ZWkGMNGu2aUrgQ9m
pZS/Wb5UzhfLCKVuCXxDiYjBPEkmkzPb8uPc2VnBKMvMzzLplbXclxbimovMefKoASX4yEeVaEeA
Sr+9OpsK1ZihZMPkDCjxU0r07vGN0xe8DIwDob8thfGRsyU4v9WBBx0/9N22TVBzfXUBlLCX9HR5
7ZXJNjshfCcVygWBuBO5GZOvL7UicY8TT5YS+7vsDId5wazQIyM/HX9WSr6+Gq+Cs5nmpbkm6B79
7txTOXbFaWSskER8t3IQ+FzozaX4kJZdkD6mSidRh5fU6leukJ70qg3n0lO7lhJoh1VXuceMCCwG
O+L8ofyA9vqr5nDlQ8GNAcQymow0TqvgpyA3y4ISgDXKbd94T3/7mb0kVlTxEcEG0bU3s7O94FpI
UUmP1wTObMHtBasCIPKbBN+FaQwsMxU5yKe6k7M8NxiMTPmsBmcaOSIGM5edRFOAYsPfX8bpwflt
vFTlW/CDTu/gnhQpNZPfgPX+N/EgLn8GR6y/KVSioG4PR4HUw1qdlewzTIYOfiZZYdTJNSRqGExU
jem/jjHxBaNmgWsZWsK1xvCqxqODqT7af9B6V8Jj7Pey9/YOUFMVudfsg2k6xvpv26J+EyH0mMhf
CY1gpw7UlbDLRmazbu/6lG7mLWpdu9SCLjlKuGXdPIIqHQg3iU77hsTWqVZuxauFI4oT2X4hTFAg
yuNsk+EBbRNHxriw4lceMITluJ6T9ANYkvKdKNJDz54xsyq0V3CRF4eBYRYh6X8k9+xKDs8QpXfy
wl6AjuSYPOcO4hamVBtanNn5tWnM0kFZdot8VFmag1RLtiDWvkYbJ7JUbkAdx/sE9RSnA9T7QGXX
DzYkvNi9fb15EsKyX/d/iVVKQe2U6n8sYGSXaebW3EQsXkBuD5CurbkBfARQoy/WEI0tVcqU58v9
k63rVZdYu8LXvsi90GNKRX3k1Gybml9Fh0QEDyWlUE/Rr1q7dvgdHzdqMZP0AIoxDxjnmuNyj7s4
XKH2NbD1LWVqFMI6uaaDYqbLIsnbp6eBABVL9lpPRPx5DB9jux3hwrW4S03GtGpEh4Z7KdK9KXOj
zwEI33hVWQiPE8KT0EItJ8U/uXFJm7eR0jifOajmBg5uOpurwgNSrXTOlX5F7vl2EzR7JWCop3NQ
f6QB8c1I+j7RAZhZJ1+f85axNEAdKreet3q9WfsDI98JPeFv9eORQUVGShKzLbFqxxAYu54OuJY4
Vl4lkXZRj9XNUUFdc0HerAJOE2bV5q2Io5TPcN6PQL2EmK85nMOlhxQMt2SPLA+BskcqYMc43MN8
wuSTsOdAp7LGoB24td0FDqvtk7pNsWL9Nw6tbR76NpCjSJOs+JXR2Fw8sEnfL+9gPx4Lg6c+VQct
xQblnSQa/M/jQhH0yfJZVafoupqyP02EaigYwFfH/QXbB+uxNxx4VAsUspIXqKuWu9hCc50mxOGV
ERERdZHQqgYTKbdy127cY4ZPLugNie7bYhbaO6IWTkCTQzgVQuxmhDDQ4K9c20+4h+cBP4rISCzS
NY73b4WWG2SpqEwEWlK403UnC5lK2uuWvQl2WSBQwnkTFTCpkymJ4FwMKCag54fokbGyH6R1YIZb
TIpzQSJXk5IZT0Yn8dT47qE8omsLl5Up6I2Ury5JaioMgq68MXCV2/T9yvSWe/745wbhwXt9Yl0w
QsBauRSwB1TQ7ZvUc39h97HMaiIrtgJyTwsQzQmPLLR/WCrwBX3XKzpcid3zWTH2E9eYM1hSrU1C
EchcWgxg2oT8ysy6X3GzzwBaWc0J/bndJBpeD1L51AijdthOYZSEsUM+AShHW0daDh2nbvRUKNQu
+KSDn8fAB8cT+/E1h9kGc9fkoF3L+3T0RE1dZkIlMwDLM91pG0AC1UfEIR8w9Tf6L9+TIf2vTnSB
/awlzZTlqv5Ov1JxzFYM6vH5baBw7ooJ3GNGRvUVbcOuR0YzrlpRr2U9hl+4K+1qVFyHDKbF/WNh
09YSvH+pk53u7lSHLNxKaqhkJEUV1TI8BtzdkanYFUPc6fLHxT3Nr2uNdR8VI9VqXmhoGR8ToeSY
PhFR/I6pW7nFJFAV2eXPphsw6CiwUTudnX7DcmA1pLlcIhEXfcOHwbHDitcuku71D63nsZ++r7QZ
NgSQgSX6Nan8JP2RhixnHWAjkCmz0+IagxXYgei2vicAGdNHa+5c+KR4fdlag3w3bPayjRCDhaeD
oDzmjaKIeKv+MXNKAAMcCTmkwwz07tjh+QPs30DD4gbAf3/V37I4msBjsMb68rhb3x0Xy3MkWR5f
4xJWSrfNVi/wsV7BFVbMx/JjYAPQU2TY4KRKvjfJFz6zzsAgWvTzSavs16H+16JzEGUZRlLwM3v1
MAIZEvl1AX4C0Sb38hE5fvFmZ4lPIDErwzE1IMb5cAlOJxvrqTePJS7jrjqbFuU8exoOaPbfYjZz
SNMHW0vPBWEGVna05op0fq+Vsa6lYw3MLKkn1X6oJdilgGJwy2nfvjeElbFaVpPc21OiT3o6g+1U
r/3uN8FEwyMLhx9CkrvOzm8AMwqEDGJeBWt7++4SioeGFcuUtNcGVUgxGaI8WeWf7In6fN0LJc9f
qb9FeF6OiJqOl7l++YBFsu17VtGoOKbwAbr0nMzZj2aU6pzZZaBSMBHzD5L7ZBM9ieREtV5Pf1kB
L0REB3Inzs/K4m4w6dikT5r3ksnkn7UpDWHoVmiwL7MHkZPVf+wG/qAgxSnNcpudf6KnSw9hbR0G
55X6ReN4pQOLOf2LiCoYCTRlWWB+XvKeShcVhfPz5XmzKae6Js5wtSax/nMReIJTNMBwPf7WXoAX
jFbId3F3cLlrCE2boz7esfG4GN0QrEvrcG/K04/f++ENXXQ9fZ8/eN3SIMIDJTEayPrSdfKgR/WL
5CgH+a6m7d0+/zZMSKXvdiT3JXMxacchBwrcJXEcvfmbYawX9CJw9HTpcGsHgM5IJ3nH77srIJXS
Zq+pcI1priS7q0m+YWM4ItNDsumrpCEGF3qZ6XSQgCigqsEg5iE5bj6v6WNrY2fBFes7DSxXuxDJ
MqFiH5bpK9E45Aixvnyq2cLtPkXkwubbGlPUGHrBSfW6CiPyfVPszMbhnYjL2m3qL1tswh2bJUEP
1/Um2wqRH+NZh69WpImuHbukz6i3rOOwSZ9TUUSkYRxJpW4HJAuZlJk60MO8qHy/wsRGdiv5EuAg
OQI3pLVTvY4zI82N4JyMi8GFE+azX+2DMEJ5+stGqdUjeX810SeF4eL1djg3ZJQN9TD8aRJPW7GG
dJe3XlpVLEII3dylARG29va1Qrv720PyEg9tmqWLPHbhiT4nZdhFHar45GT4E6Fgbb2qdDsge3tb
88t9TORHARk1vtoOK65PfEZaqX0vDUgESBvFbdQxYQzjyu7lbg+XZugE4AmZxyGIGPIWke/VxueH
zs//OSmPfxjkVZZtPVt72EzhQF60xCt4PKlxvt0lUvCF0PhWCaS2ASdNV7cwzGE3bWMnaeGZtuNE
0nWiKGIwTimjC8ufEjGH0g9CigHkVLHJ9KMe7zaZ2+z9rSdY0WXa3JwztL6RFWW1aHS9LxlwMYoI
XmxzMLUChNq+EwVrGsdS2ql4ZyRwjkSdDQSHvASCpz91qmmacYulfHaTe1mDNLtzX5ooCagIRKDC
oESyRsG78wuNhKd2TUNbhgW60Uyi3HtXYJiLNuol04C+bph+AlCY0Tt6ph7orkXs9cxeBhdU3fOT
ecITKoqmcx0j8kiQxiWPFPhRrFomTVnCGKYRvuylSfu4Qimf6PrBYi5MW9RIUzzI0dmr6V8pW5zG
Wy5qOPu1yc2E9OEKnXHp08lZlake+V8PT1+oUH20UnousCfwpjVlTUfTWIZFrKG1lBpSEmfoeTvD
75pAQNrO+N0mVPU/sQ0CgHaaN2BqhsUJIO3eI9CJm8nB0iWRACVODqhn0XPIQgF5FJYVQVZmLImx
8kU7EbXu3yXDrsMzDfRnxuhScB8SRNjqPO3HPSlWBiSZQSwTbkFxpYPqkzOwsgC50IOT+XtGnaue
CTQbHwcSKJzt8qsiEU11MfpbHBorlXW/lgZb57bLD+rxKvtxCNjpj2wKStyw2S/mHAGgkgvgrfPh
AVdXUtPUm6OdCqJXeSZenoUdcwYpwzpHam/8k+i8pZLdhT7xb+F6CFljG0z0ZN3Xe4ZOG3k1ToQO
3Ylwti7TTe5RbA7XnPnTT3D08ts4TToCeTDr9s6K2JajObyG/+baSS2bFypoBa+A83OAlXVf8fTm
QDE6sskjtzFcBPSW1F3wSAVNXyHetwpPA6+R75Rx/cy1owOj5b/zE84uOjchbRtC8chbp/PQ8BpV
ZtE8rnCsP+flyOuHndGEB0jn3wJp5/e+nTXgTLp/4sKZq+39PjSt1G8LLFeDaPI2kPLhhFeCnGmc
gsDNUO6I5ezrvrwzu81vNc9yNScyqNRLsGL5gxx1mITwsWydbRhR9qzPJcWWTI3kxgyetYP7XcfG
c9AjmZILwxKqa84rMOAYoPzH5RuSGffFQ4Xu1FKrbOc/RrPAR1ViFpZyHWqDRzWBXthVJZPv5I3+
uaOweaVDpSEkg6bmZn7BGzdEu1C6q86DBYoSRkAh9oYLNBggKfFrOt1p4xS7eoGYiROSKVDC++hv
QTPEdgABJScdOd4UvLMPPno7FYd3ppmZomDjeVAWCK9EQWIP6NHYre0f5s7wJyDKf6qVkmBnWYFT
aviYoUZK2lSw3eF2Xlgv1bY7+OT84B6qSuN1Hy8pKf0N148xh3Q/Fdwbi/Mqs2+/z52IZLBYrQgf
cr6zPZHyWo4V/cIo0KJqId40rTmS8H9LfyMyRk7hRFf58eGFXmok3F5KUmGeOvQkHwtWHWgu0ekq
V13UpQdpaiTC6VmlmxYumVA+Rrs7uRu7d28GRu4woGq5svWkWgooWKh093mDNhmGXtkmbAwmmieZ
5QogF7t3FAJXejB+pn5Tl/QMWy8cmxCopU7MF/ZlqDhunAohBZ6lbdEKX0P8HY/rfQxFT0OsX8ji
q5k8zCUTEKcb0GqJ1ZHR3XiTOdLVJAy6qkn40dtK+mZFx9KSoTHvHn5RH+6OdGtHVRn5KubdLChP
otTO/VfBcV18eV1G3gXk06kfZdfikwPKky/NnEA0cwlapIznSOMcnvCAp1F51D/pjBCcLZwPKk8E
gbhRPu5nB24A0gIvhTdPsBZEjiDtx/VpFSWhlRd0hfbSl+K/W1y8TjEdzRx5Gx+RHNX+ZHaegCIm
1gQ83+l79pfDifbDka87K8fic3FiU3cYd86K3pQZgOM5BOv9WjBE8JJDiVytCknZGeM4mn3kvlV/
vVx38c5w+LJm0JsFHB5tecRtYF3CIFaKPptKHCsSRkXe2tZTzjk78EKnUBGJ5c5vOzgmmTEm9jkp
TcUXnBT2q/RF7KdhT4tBCCKh4qyxTeOHEPf7yaEsfPrFmkXBY3hI9EPUI4+n6dGDqNVphp/PWRol
rVYo7hROv71rNzItTBimnPSh+2pz0HmDEp7vl72ZR1BCetErBmMP/Fx78YZrOBn3J9yRTdCfRoMX
6ia2+BOKFuea9PcRNARys/BHrZ8PyCDdIO1YpHkFWBYIbmqNZ7Av3kU1W56w8l6nJ5sB3KAxn95G
9+hyObPVZf6dCnDZgb0XZ9xkGKH4WGQU1+ZOBzGVl/vToiDMBchAj53YNM5sk5OyCU7MU8InhWK5
sYiTzoynrSlb7r7zRZdeUY7Z7wZAX1WfhFawPNOogMQmUrYtpks1y44y7/zOJmb35t820lgyW2KE
6UpEySPicqg68SNCqjFZbSAxToweGWZN+BeYSKGaavrAUjGrl17HaFDRpCvu5JSSnKbcYVj+ayXr
sDEXKo4b1wY7aIpAgA52wFa1R3QSj7dOVDeKQxwNgRC/Hsi80NpLmWP9FpwQi/me4FpIP/0/MUAf
kwEOlIIHj74RjxXcOx26IpM+q1/Hu/NFqtSmkp+9ntPe5JO9aSKKiAG1W5OFCpYElXv9wysrZOk9
4HzcF0Mz6E4PHNojaKwrUWovHmdioas89bPws7wNkioB+l5hziCfez2IpvopzOg/Yss8OJv2kWzI
R8ncXRlJU66IYjJOpfzsq94eHPNncXY2fATQ7iJO7TG7tLQ7EBNwBoL+UcKjwO5wmL94dLLOVNya
Pt6OQNjVjgfiNSzPnuhBuIsKIk2tBwiNqyQV8XZgibEjjzmhcETFJiA8zy6a4eN2BBrvUKt7bjll
26OyOWdW2kce+Y4VOjpNAkc9cU0ficbDbzL+sAqsMR4qtiSP6PDnngC2PjtQk6RU4gIsiQx5uQiT
aimGaUzeHDZXKgrdptwK2VkLYkFBQdqekKHmHwJo9YAqD5RyO1EgFNRVGqZNt7yCurqsy2XUAp+6
bFYOCqTi0fMSH4vk9plaSl6wh0pzGjFq8LW5KcMkiruCKyEJ3+G6TzafYSGjD8AfAekvFPWG0wSZ
/mXTXxSU2qE80XYrSGa2tCRzgnb8VmHKGjAeATXl8lGu4RC6dD7tnhA5/Lk7P7g2xBBh7JaqCdbZ
BnPYCHbFj4tUuLvw7hzLPfDsNE7Lg3dh2xB/LYmfNZNLNYoORgVjsdewC3pjo3j39rcRp3I/40Tm
t4wv6m8dyc6aH3YWdy10o2RTjSEQU8EfuSJ4spdw9vVT5jL/b7k3j/9j5BssFUzNgBbu+GhRDQ8M
/viHmk4YsLalt7a+TOJtevnbhimY7q4Wb1nrDMHBo42brKaFABIpA2a9/U5OxSmWr3Jp7DlFOK87
xxeLk2pagthQF/sopOtBPX12jFUHkoJpMwAaIaXTFLddv+CBGR4DdfJU+tdv9qMDdTc7sxOZcwW8
/xkF9252wdGjbqSZpkGNpd3nLrgmbClRz0ed0n51vO6PZh1WBvkWIc7HSilGYYowNI37uhbKzDdH
7Li54fYC6Bm77nD8O6YGWTtYQ8//kO69cX/+Y9UvsZ+9NNnQv0GaNysE7n+SeX5vXodC+1wSU7MJ
xxvav5QT1v5gfSGG9DzhvZp1dv2+n37KavwkImCNTuitrze9OAJ2ozrv5xa/iJxqZ0YjCqgFG4bQ
u7Ag6Jli3kSBVpxayNlh7hVkD2pgzWfldNn/zZHF1SAqHkjfpqIoPMIC1bl7xwG7LbPBFhOHOoS/
oUeWJDCdBtwGcd6PkLcNCEfXff+0zQx3ummGsttRLOS/MgQcS2/85lA7pzX1QHBIzT2V+0PUEOtp
oq3lk7TBTsx35uSf+gu+f/sYN9Uiza2ZmkTuxyPJolw5cAnKKZQkTT5Re17TxxFjKGE8/WcA10bA
q4ByjrCGQeYqS/vteHXsN7qW7OdxtW6ivL6v6D/eJgvhrLzWdRXtsgEoYenJ55X/t5Y+9Pdf3VG/
o6ySIo5mRX/glMukdFS+Af42nK37wryquGwNGiTQ7K/bFIckGPrI59MszCu3Ty8sHOhdvL5EM39e
uS9JfvkxMtQ6xsrv1tcFpO5U5FQbTpL0lTclwARtdwwcX77Xl4UJytxkTDnJcK14ZMpoigK/AGyf
JX7TBECI2zjB6qu+4di2FDh/bqMluORAr39T+was29OkNx6JkcFexYxPsxOSjynzbCktrH/Qp/vT
q6RAs2j8nAsXtiqRKcz61W/IRLO+mwttomACKao5hXwvp8Az492gnfduSqusFbt0bEbgXbI7GyWG
nttpeI8nnEEegLhBuyFvaYq/pQKeZYzdYaYqewqdOmtetdMabGuU6zpTSysQCcHjq2vVxp6Wzfa/
kuApbtxRQQirsQaGXw+FZAyfQWxKUHgIP5uUaIaiBYEjWjqF+20qVUeZrVnPDatlhWqPsoqjLEug
Mwi8wYW+p40YgfSq7DNBm3wQ/K2m6CWkJvKkWqmLTxOISXZATdDm3Cg6cLo2vKAGn19Pzr5cuon+
x414qc/EIdUSBd9PjzpqKnjChztxrqleszIfuRL6vFGaQ6nwnLa2FLLYCjY3fwC1X5iIopdywqrr
8fRpzl9gdgtiYZT4oxScVbzWFRDtwtbsaUf0lgThPtso1iEy5U+Fb6k4C9mlO7r4sb/GVY1mtWB/
Go9PDVxNOb4KwKVVb2lQMULbG+LeRFr720v+XLD6Qkncw2jlWRphvZUITbIWxMsNpgTcvOxT7bhy
shcmiIAm60cSlCzRmX1nJZ1k7dsEoP3ZzPivdkXND+liCawqmVVg9CAS73qP/YJ5nMYFdM0YdHBk
6R/t0VRWZCTDGZiMHgY5c3pp3e8VTPWiSC8OgoZtXoqufVyA4RmBwXQjozoTkjMvist1akcnk+Xq
9vgljLeOtof3Dq5ialGYBXWx4yrk0aZcatiYkd2ITgRsDS7H//k6+x8MR8zWoPlNIx0zfnx/c+H9
XK2CGO0PFOLvM9VwIVvHPGve8k3WmPMTAwGxg4mhwmYWGlniTxZwBZOUujdoOXKeYnemLaQ68N1C
Umz3TSmvXGTIcw7PV25SYCkjANQweAlcs8Bx/ocVTdD7LyW87AuzQ+eGms+7dh41CCXlnLnYwpUe
cGuFXuBagdyDhZYGe7fqYrMN/V5ldLClOy4+uaI3XZz3yEZc17NUfO6CYFyGTpJI47cS8IxNk2d2
qMnLUhfNN1edAgvCtviyXDy6x8XfDuAzdxY/ieaAfLwzmY5h7uLZEKsjs2U2vQGN1N3S8I4+o3H4
YazBshonqrtT3aT3OJ7llHnDumR1tsjkGxVuXNbWgTP4ZgQARoyYnd8P449PF93TOrFA26MnYxkQ
iFbHsi0NUiN1htblMN7f/DJOzI2ZfGfzfGpp/dv/lZb0Xm3Vdrd8bQ33nCtbPgMsl7NQ3Xnci2pN
kGRexEWHfYYb02LGle1ORYmszVCJ04+TTNd1XcUQUDrVogU1nwkpZpbeWSdkky5gxkmwWEEp4zMx
aGj/db4g8pwhtEQX1a+bRWicd0/CGarfw6aEj6rCGQlAxQ2JnaMXa1acz3yFTK3PImpV/8Z6wALV
2ZP0UWvb1aoTXtI/ZLUwFDHORBCbvfJYZKN1hy8EtdDp8EwfvdQpxuOB7HiMulSAjVIMlDXYztQ7
Oi4GxwotvqHNMrppWFClremhJPGI45ireZbJuJhHmdUKiL1Kk0BHaqa1kVNlXsIkcnIwIplipYZo
uNQOGtRXukzXaF5H+GJEEHPraaGZBlBlFHhTHS5zkoo+PBhlHvX78pd2TGunbwdwTxEWfpsbQ8+U
b82ds90RIMR9F/Qr8qDDswnzkILFZ3ChkYnIZsFoM8T65X5HgTjHIRGru6Hq7jUribKxoaCaqHJ5
MWBnjRvINNh9BVRdPMzqm+yrJIyHH4Fg/juGQ7BaXjQvNgMKko5O+uk/3hOinnVqagGnWQIQemNk
Bs/P6dfaGXFmBKj4QPU60rbSB3Gjh+Kv0z+KEwmGyn5VuL6yohhXMrxrCbCr7qTkQIV3iI8lsML7
zk2yMkH4RLoFcnFf1cVbdZuHoDt3Xn1g9VaLYaEUtTDPg6oksZjhDtJkeZ4yFai2iEgi5eF2bhFX
WT7VPb2jqGBNfe//4zenyhAot/+eh6BCCnd51fkPVnjfbNh/rWH4+PWqzyFUVdaSBWPdGamcIUtC
woMK7yd5P976xCQCTuzINEHTXWTUaBCH/QBlo2GBRsab5Yg+JiJnXfrztRv3I/wuhlaaSw8AS9U0
ZGfr7YN7u/eRO63eI2YjaEWrvYogEl8PZOIQM18vWd1HgBI56JNOjGzBs16I+LfxoLLov0+f76Uf
ck1Uj48wKMfzejTUS8HWTPIn5U2bCT8poDQwTcdK5SPDNI0Mzl8LR8vH8Y3qKEZeACA5mTTOAlaO
sU3p13ELJNw9Po5fc17wc6zcg1GKZw3P2xnwxYjv08um4aIjwds4zlnNjaMNDLnXAzXhZQTpXK6m
QCchaAdaw6kNsBu0CRC09TXmqASAffbUgJCJI/CelrCjQM5pK2x88f33kTGNzF/+EhS01CSUucGP
WtSwa8/1FU6WLHWL5GhmgyL+SBnAaOcxuRvVq1XHLUQWKGrHEXb/x3rqQCjnyWxfL+9uNAKAWbsc
WVal9U5q5G8ExbQHmXNhSm/iHnXBjIQBTt+zCgr17bg+8eSP3r9j6Vh2ZmCc0WDyN7aKdLvsBi18
Z5bEmWA0W+ZHNoyMLrZawGSTBwPJb02LFNuM0NtstrUyHbuh1xFDEsCmoiYpEYpha9aWsJDRKjuw
MhllNk4CdXMRiggfpIz5sr+sfqAUCulIT2+ikN+CzhtTjBxupO+Dy2BmvVJgH42PD6A7Gn1lMtmj
XESYCVtkVVvD7sBGUCyFbHdiSncrfKQDrPVip9v4i57hhtVvXr2sicVrDciDQEavvlpOEE8VEuMn
7YbNgUQq8aMOPiM8b6CL/+YcjHePY5TT69Cc7Z+V2A7mBRxx4buntmChwjVhShnvjRiPKBWT9YtG
GJrsdq69/lpZNwgkTzRDaUfuAf4+Gxb5vIoY/55OHxVTZwI4Wbyw+qEY5Ttehm76dwUAmRVahZRT
7X+mKFsBkeM0OEpp2XJGcepNeJv2gJxsmRETV0bIKsyNYhAwB0QANjpomcQMeaKHmJyAwbyTP0Xn
Nah6eaEBuKKOgzdW5TeA89WLZfh7DTHNQeBGWmif1bkgXT13pNvThn8rz3ZgBnxECpN5jPKQasol
RU4fCTTF1P47PIeab2Hiw+0fc7WB8CyKnsfgs/8qQVrbrLf01wA+Jp5tCdHHRvuc5XVUT0WPfWzs
eL1WrmHGaPO/eZwcJ54aaWPzV49c8AnKPjQtZdxoij+chjV/6u7jXmukF1tM2rVLOjQaJBoSeOrz
FK+gQGz00eTt4Da8SMBPOOQkjXWJZGBPWSJjczCWzNNa01v2HJ3aXfH5xLQ2TtJQmtIEid0DdRz3
xqYtDLhVNXc7bOPwk4UBkQi6sjE/Lao3BZa4AG9KNUf9Ib0+RHWqymGXH8XBXeKOn8N3qaM+oLX+
u2qegv6xrliadLr8WMKf3OMBJsP9EG+CnOMxQedu27MbPyGwpLoDsZRmiX4YlwJsNvj8ddQLWvd7
cAl5fWzB0UyrF76il1ku4dRAKQw8vrCZf/TABX8ZNfEbRDfuSwd2lNG+MaMT3swevjk4ksjt7Pn5
K73/Fe2LA3PBGmTDXDnVeZ7qG7BCRifhVXR2wZm6E/oUevxyVx+eARGqxOTVM0s955iQD03VvMtw
5No1N0TeZ7zIcJJWOenMH5Ma4K3jGrwHvWMT+U0NLiuvRJLLwCKGp/7cz/B7+KJ4H/6J7ExA9Nvp
P2tyBsRoCVIbCQiueXtBCxAN3kCLZMkHFbjnexqzgY2hqw02Qo0Bj18ms9Bpkx+EVfGpMy6xCzmg
JREfWe9RIPyyB271hyWWYfnhad18oTc4sgWwYZiTmrcjhD+LDVdan8k+SgK+YyigRdYx4xXa3P+w
200iBLRCJyHo43Klc0Tc0K+MPkDZLTWUOyQwq3NXb+fCdOai9pzA9s0LTeqMfb6MtoBjyIRdaxV+
v1wr7j9tiSXdp8AURFCWkWC+AExXHZw3LOD6KVzLrAmA+yIIHnWqVfSet92kvvPrzBOnSulI4tj1
ZV9j7ZXP0sff18cziPCdvBK9NY02s/6hXoMJKGvpJlnFIYr7OAHy0NqG9U2awpZZtEma3YKu1QF3
BkQpsuPQmrad4ugrrrziiDiBzFK0e55JTMQJhTUYhiPaGjWRk6Xoci28xfCzdJXjAlSxc8PTIsnL
M2rW3leIWk7u/1zo5n8jEUV4PYgpJdsEH/v8FMcur94aYM+hH5Qck9lrsRbZew/+A/MGVEuaPnAY
bjN+40rI1oFg5CEqZmAtWNMr6t3HTHMjpxdg1rpG9uqEEupx1wtb3a8KoLmAATxMCmW/Z9Dd29op
v3q0taIj7eA7zxy+UAxH237OZGQuMTlaHBTynWyNWHoLij8qqQsJ/Wz/8cEEaJtNOVegBlbsppYI
+SqCIsUYOHVxJ+Io9PaVm1gXjj47FdnToClDhfY3EhpB6+adtWrRnTdC05hrl7zw8/Y17Q1JF7Ep
acTemcjen/ouFru4qeeLk9wn79hq1bGra9gkb6ccnBoEvhsyy9m2lhFm7vZnlbgV4zutFqgOozLM
mYRZ8LA20ZJCqCdk5ENeAKCa29bFNIg+OSKs9EHux/HnIMPcUcvwbygLaYOj63uxBw/iXvY8PwQh
yy+HoIu3cWrJyfMwSjkpzQLzM0f44jQS96m39dBXtJEsFFfWTVJ95Xs0S3NrrMWAFM6XMBq9l6In
Pwc9IJLnfNEJ0pYPO74ST2tefXQKPPFumMq3JVd3WUkC/5wCeA+0gLHzAhXnC9c1R/Y1AB605g/Y
LgXxKBgVlPKVyuiZe/mzzHkuGtUAUs/RT6lH8wvxk9nwvgBcOaSjS8aHv4/6hwVDf9cbPGRJiqU4
CuzLf1VfdzH3dKClP/mHiRye5uDTX7nBWl8oHCoUd6UL0zHjs7T1Gec2Si2Aq4SZpVOexkPWPzKC
tkjFiwnpVozHxXE1pN8I17K+HuaOcKWchL+t2q15qZrZTKqgzV7lQ65nNnJz8Hp6us2qul3fdW/7
ofXyBHdWGa38jPzz4/xcpsDbRodIHBTMkXVN0ORY/lZ6a0T6yLFp0dLMK5kc6ySiB0AD66qcU3N4
yuUWRWgNR51d88eKDKeEFxzLmCw5s43EgEFelcjtX5sk3bFdc0rbIPhztKw10le1TVR/herz4nre
B59N+c1JEHoPIJbjlBZYpwcHSquHIlteBcIvB4wsHYqt9QTJQRDDnHoGaDwZ5Ebrqb/9k83n9GVY
8Oo/hFK3VxfKi4j5uGWeCRj+pXaSrTB3ezSwukKIWmX+HimLpZWR7F4eYZBskSh6UwaKP8PqLutG
tB4OPmCWeY+FGsidakwv1UuoiU9URHhUINyBN1MdL5oJlHXWG+YoDdVaE+ot1O8fU6TIJIC7s9uI
TCUYAwimVghf6iFq2EVhbTNr2Zu9jWKdI1KZuidRAU3ZO0KTjelE+++gjj+uCOmqP2uWibb9SKBO
0ApF0x4mDNyhNYUkCNe0qSX579ojIHG8tWNzf2BI1Vb2PToz5eu/q/Al+snqfNfCzzDBvJlFB7Ls
J4cn3zZfYwJTkyNUPx0i6t/zljUxO7asp12ry0XlckcTG+kjB4zwKD8en9JketqhkZ52atsPmlU4
4IqXvt5eyI5F4J+BkO6dWR6rwNixWWC2+ToifQih10FB736rT8E/EPNYNu1/QCNU73vCXWgFLa2t
4wY54fzya12abZmDsOhhesLBC3au/1PRuhBvyrRVbW/PTCoSGFxG8zc5DULsXLvGpew7d4pY2jYA
OwRWf6BYSS0qwMI1f0wByadoMcq+NFU8ptZAO7iBaHOC7S0Yw51slUmm1+hgzH1bBaJRUTPQlwVQ
9Rn+2Szukn1nLnUev1yydECUj2jT7zvl5PFNIlL5ULgRho/klNS+RdllQautPQEV636OZl24/rUH
5KMP5Da1HGHe5DzkfqolFlVKQHmoZ5bY2OFP4mmTZqN7h7LsJuUNlsraOWUZDdzJcSiC8Lz2hhpW
1WtEbp9hR9GuvF8N1d+/6cftVOoAR5+5d1njCG7OMns8YGHwmXs4He8gZ75NraYz4yN99Z+IT8Ky
EhdPfJnp4T4dk4d+qIIm7tunkYRNnfbzaQhmubL6eqspXaak2H7JoHkJHolN3LsJs4/UzLrc17MP
K23u+ruq0GHFrUP8VlsY1N87RayMW3mtTqbHdK5XtBiFfDPnqJquvc92EHY5J7ZDhgvVdggy+m8p
VM4ACQjQmM6eyPG3pfurk9rQAceVBY6N8A8CIwJZZobMyxjijrTFRS/vvAZlZXU6K0DnIaRT7arO
LgmrDbnZIs/MMj+xaOsmgZycGa++CccShBWmTATShmDwZws6CcklqXMlwa+RQmgNOjXMC/3SiXG5
17nfi5nqqyEvOPAsX+PyVFBthr2OikYdoG63MZq7TFUvsEK9IeJbt5JxgdFrrdgagC7jyUNYaB1J
xdlDRO0yn7UGbQTGgADBWHCRT5RsOb6a128ADfLLmSsb/8vlebjveyB5QW6F5zrvnaWkdBb2Qeo2
mYcypJ5NUBX7kOC7aQdWRHrNiqKJJYJhFZfBWtAL0PJiGr5VpN/g7AUPV1sU6KxqOCmYz7f7TKEC
bZK1jproiRD6mWT02GD90yNgRpGnT41IMCSzWXpBrKfiqL1kFk/H8AycpD5HkucVntxt5/Gr69ZX
hkcAtwN1Gz0Oy9Okad80RPAIphnAMQr7K2HfoUbeWCseNxBqSnPaTc1bW9FzsunRYVoEV6BAHtW+
E18vNsNJJqHr4o49ivYy0pFbkMkNolDrCt5VM4akxcvIimXXbm0+DtW348ibUaejGkuxQmKfQ5oD
wD27rDdNxYJiZI4AoZEyMQ0H/rVLe1THpheEHAYCChhhKnZAKxCkqo/yDGl5S74wuFykgoJqeN3R
VJALnMMusHXcVCpV4lGGkoU14YEFqikilFH6a4ll70N5eSl8USTvRggQa3LbdOKifzAVSXVOJKPH
22wdTf9b8IagAVLUPBaECQ99Q/7Q6lEhL2sKLPRr2hqXJLIYHJaRb9glfAwSU0wI5cwS/DSx7p4W
SHX+Cb8Qjd2g5rEF8YE3HUiKftVMwVNbnefycDtIq7oHgHCYgIb2BkjklFUS7XCSgCoO9IPDb4Le
+EdgrIDc4PlCex0AiMATSlnmOdn0xNrsPQf2hNSwXeB3ucsixi6LyHAvsugtYRlRzeHtpcGua89T
I8vmp84CGdeVgX++ggxY2Ish5hVTEArSae9nM2r26tig2yQYafGxyWB0/NvixP51Jri1OVHK+QU5
+M1WV11O4NSdczigt8VB+TY62eozNYo2sUctOBjBI0uKWWOHi5z8kg4yL8AgCCo86WJ9vs67mrIe
k5iaAEOtXjVqdBL7B4jV+puwPXbBWn5Z00sjGwyKTihKX9ncY2Cq8OKj3x4DUdiTXKumqnjd7Vmd
FQwL9wb/7HeZjT9ZWNF2iAClM0MK9A8cvF/VhWg5KPaxBnSuQi1SGaPUbdxlx+UkVKW/BgZ44Ex6
+s70TJSodmrpPbku5D8mfPV50y8GZiIe/y3eNdbPiPeoAAFw2qSTBvTvvSzh25x0KFrF7x/+5oMi
hhFbWVHuaowIMtOYWUmhPk8dAGdqU/ry7mSh5gB8H9JemtVx6xyUDHYZisbQRD270DCAJu61aoX8
hlknDBv8Lnz9ienh7RTZ+yzy1hI30S0q6lLfHs8YmVXTruMw6ObDVoWYVe9ckgI1qfzpgfhiGPOo
BjDsIogYdkiRdWwOaOk83EdLJzQ2d+YsJ25fDmH+Ry77cU2t4L7aaRQlOM4Mjav/SI/55iEhtVgi
rJyeoYwXyAFqqAsqCRcsjB1+1rlh/bFsJCEQzgN1KlZDzgP6/7WVaFSD/kggEfeJaYWuQq3e9KLw
BZYAGDvXx6hoDVE2VZNByZ2upx/CdteGbwob20nuXTQYfY+MTnU5CP683gsnG6Fu9hhAZURo25jd
dS8AZS0HSUbZ7VVKmawyitNmKuiUf/3/6Nsb8mqR84llidOIsqKFPvhHLKtLc7K15kbUaNitjUY7
2ekr47lyW62XLxvaCOk04+gETP7fVG3o/uecGIXPDXRCxDkxf+ZKpLOjj85I3o1k/9PkYKvFa0eA
Z/qoxmn6NDL2HdmzU5Xw0l9Fh7fSiiGgJCeB9F18eb2lDUJYy2y8cTLHx2xkuhDEE5mQCGezJo5I
0UxhzIjiqkb6VAKJ+b6hhmKTISdOqmiYnFdf18pFVag0LOGvpbYiQBPiniOpeiDF4HthqhtXyJhk
Mei37oksYrKRQ21RuRdEs7AeWWU7rqHpc77L/eP1axRyhUnNuT4UmNcXRXuJCUrJSggSW2xkXzZx
QgIg4i/AtKb8zdwuiVzPmuSLoWa6l9EUZNcVTPDRvKKCn8yAoGBnn50LEGdOBrMoi5H7YwHOc970
OoqRDNh4khLFjyhxgJbG9Ku4lZIzeXSiB7Ygrh4x1w8iVk2SJcnCBFMuJd96mUPmpg7GMffJoIba
1xZ3IDdIsa5cqRL9YAF221MN4VzI613q9vGwkfqr71QGERMxagqFIhaYA0gSaEYCn5AePqinCRZv
xUPzKCyCkNzlBHkHkxTR9HEMpmHBzd1ozYmnWB4D0FdDZBoF3BvhNHkL4A0EB/GC8PNJ7/WDDs30
Vta7au4MStu0mnShYvfKVaAzEK8j2cl9dD17ofyxGJLxJeA6k4TZx9k+xTiWYmgudloFvJ0TE/6E
idqcbfvbF4LARcIoeyzrpeyCdA5fGbN37yce/nnGSxcSgTCyyB1uPWnPWrwy57pa43GgjB54XmYX
AUecZ6hiGdIPye1URUh97b0LvSFUo6QW1Z0qI5MvFmVoU63hA3Am8LgpHa/kLCfsfueMVciDpZxb
F8kwrXSjq0NYiDSmf0wPcpD7D8w0j/UZ9UwMUzk9cH1imVqJG2rx+Es88xh76YxXrp0AT/C0Wv/7
/a5n+e9mIdZogtspYtI++u7yeRXTbnYignFQ1lZcponHGClXmp5A3xyhDX62seJTc54bo1B8X1h5
Xy0K/jaaSFGFQj/gd789iBBOS5PGbr+wTxfJPoIlPElLJ512hdY7AhHmKGrvVqJICK5m32phzWIy
N4IIgYPnNfwVvBJQsfJftXr0YjuVN9w3RD4qSxs2tmvdHwZH1IBu2LjWxojAOg1TDYYw2npQXawE
eVcLbsKc3adl1uKicvnwROIUKMTJ17haq4USbPKlJGyBBt2DLdFC/QuErzSNg0Kgv2fCnnl56VGY
UP4YnXTk9KOIntX7LNalabSgWja+jvj0GVqyAQ4YfYWr4IMXX25KmmbAFGRdZqZwUhZip7+VhLoJ
sNGOwWhEcr6g5nuussXZ3EvnHsQZqZjFS4l9DvPHXwahk0bwWWgR5DJxdLHJ4QNMNEYMO6NsXfet
VAmkZ7GiRCvA1Ss9YF7aJjFzzu3Usm6nRzGIxfzj9TXRsXHh8j6d+uLyQeHjV2fd4RnKstgupRX9
KfiWJTw96DhIuV9DZFsal8SWHjxTwKr3Dh5qyEJam+vzqXC/YpxUXJA51s3/AK2Dz4Eyq1iuv6kx
WRWQBZnk3kvm23ty5pAHqDLSLKWEBTPLvRNvVNUgA5S1B7jwBTThvxeTsrxonGzlh6H2v7BC/Eh3
zPOovpXkqIDCxza/mJ/7/9LG6A+LCdTmB6cdwLie46U8lHf7eqYsXof7l9ODLucFq60/3dnIsJqd
YXGfEpYRYtI0IqryaQXd+HAo8mxexol/W/x6E4wteWlkf2VYMhggarZNc1ePto26Ajq7bj2f8IW5
Bl7pRAnY1rPiwtzN+iNw607bg303clbtqgsJs4b4cTPjTqq7dqjsqoNjjnNRCqNoiJogZS/wAaEe
H5wzfqRUwznLjQisGyq7cbJPc+0rLkImijKWwEiKSjjpmAkeupBZ7NssQ6jVi+mrxh3CfeHW70Nw
v0EmxgBOkL0alky1EGtzZHoydQN3FC72VtrK2UBXV3WfQdO2Q12/DbsxbIoSk9yCIlZNPWrfYPt+
xACvlPLWm181vgoG/9iiP+7Duc/imho7FkXoV49iD4iWbBPa7kzQdeSpeMrDyPvSE22lF55GlZMm
Tx9AKdsk3lirCCc+qw1jZYuhLO3FLICur8IScL6elshA5N2Vl+dL5IU9j+L30KpD2oGatfAsI/rf
VHfWtklNU+VMriu3Q1upORI56YjaSv7tuKZkFETrqLV2LWM9BKJabj6nbXzlGaNau6R1bQ4c+vMl
YznlZq8pnc2FH3RKdmzoG0L74OVE+REcMIruJWVwlG85NR4XoVBGsr/trcFMVL76yaoeIPxNESTS
LYVw9Ebdo9Fb7D2ksoTI+Zdm2qC4i3Z+CmRAV45QptmsGo5EdJhMw4PbYvkA4fimdPjwpIHDs+nW
jQQT0Jsv7HfY6LGbHQq+Wt34sD6MboXfFHzVbYTAvl6GWL4PDG9Lkut+zET3oRnEiMro+7Kwk7Q0
cctJMDNirZvw/KD2vWwUZawvi43zOU7Zi+IUIYcgkI3SSU/2L7xlYnO1ZTVxKSk8vWRZTbnKQI1D
iO179a4ftM09UBsPaIkTrZauS3Fs238jDCPu0Td14dTt+MNvO/eKz8OapRwKnJ/3lxByqPSqB7gA
KaTF2V493Mmdpd4pAqlYzpgAL0I4WvBSA2U9gaZT6gWss7SITDVyLsR0XVHZ/MaMDnI82OTbBTi0
E9D2HFTdrLL+chX5woHxRPaZLD1ERdIxMbB/MhmcdepsR4FMDAgM73KjZ/p6eOmpAcBqKruCIc9s
Uq4+xTzLf0sw2KVyQLegvYvGUH4iN6wxUuPr780In2P3U7NK5BZ4sGJqrxl/d/uwNmaA/bLHgGBl
69f/0yfSJmZe1SYpo9zBStwdqeA7VhtMObHJZimwBtPKzA2O9Y1/7UCQZeQjNFMg2SLSMZ2/U/Jn
wSvHEjzaMm/UJEcRmJ+BTnXnzNzjxJ1YCX0GhIRXiiAV/81cZ5SbQafOBvO2MnCIgDyv3t+eMHjB
/XDmBQ+CTlUGHpgV7KrLo6knlX6hO7l3j3gcSOWVZsMuqC1Lw1xxNzW8dc2WOUigASeAcmyrEMNE
Nfa9Wv0lox5t+RQKFusmC210QLM5qp10bEaGSALmbg9urw9NpShmsG8E3NtWC5/g296Xoi9D2O90
EBGj5b8cI0nRIBXbZ72YE30vTJjrt+l0HHIWyoTjsZPjAr+ohRDhQ6kREpa/dAR2/dUXw/8+oex1
wqIBfqe71lSmuy64xPz4VNXN8RdDw0vSp8AbLqC2n+cprjLDX/KlccLsdYKPvgIzLRQ90Zx5e9IY
qrEMWlv461oMDfWMwgpKSk5ga8nJ8g8csWwOI8HbzES/XXKDi0U+jwcDyKiKwVHGpwkfJz2wiAMV
BKhm/PQLHtxmVqkx2jhGb/47dlCXV50y0Ez8lXiEQCecohMGnJlHj4OHgfkufi5V8rsml/WO+Hu0
SaUo+gFdmpvpR84r6QoL9lyYhCpQPF8jDJbIi7Z15Q9klm6XAOm3tKo+r405NmYMD7WRiMHyPKXw
nZ6ENOlQu6G4UbQQTI3q3xCbSsJCFLPPioNHnAc9t/RdGqgjUntwpaVbyHOrUKXBAqarPyjHWTVi
xzKLwIhQH+DCQXPmTPkcTssyXIfJDixAlC9ZaY5Y5nw1IxCXr2N7jOtdX6bHKsL2GswSaHu0qkGf
RZZsHsq5fPEtiKPXnt2D5A0ky1ZEoUkIQb/Gd/+Qs7s2wrBuc1Ub0zR4ECdKb03Wv2hrQQd8a6ko
4UquJUaK+FPL1fKQwzt9+fQhGwa9uQ1kWILKK2F6PmhPk7CqtBbO8NhihDPqNwsBYDz3HnPAfrkm
16ypnW3J0UdQGmnmk/T15oqusF7taJq/4yqj5thm7UaW9RyN17LD+W/oRAlALjqNLZ+Rexyip+Jf
zzlQebbMI5iY3CSA7i5+cN8axazc/uI5sbiOwoEoYpZqBbwDAgjCQd+VoBT1iVVd26PVEDGhtk0F
CHemwvQ80deXVZYIFibF2hes8yCSBZNUL74hHLcDa38GOU9c88VEqqHhmRI8AAzZB3SHJaW4wR6L
wKhEC1x1xNtpvyWDfU1mHBwrXD9YTCR6OehcNjDo2rp8KvApAWiql7FUoWu18IbZbX0m3LPb1a9Z
v00xV6jrPsn0HmU5wPGqpUmhLGzHYmcEahFagLrFfadN/grASVgWOdym82HTaVaWP5fjmQx8h8MC
BWZtPps2L+bwgbm3f8RwmH7P9+MW/LSJ4KYiypC9Zbsi7aTLuKhBJvjK56A5Zz5pl0fELEJV6xdK
sFQE4ETm5yaaDD/X6B/nSLQoLT2Z1hx7/2Sa/O9RDi77fE7RexTCDJr+PGcolXgiq6qkItb/72rG
9j3NynrSxeX58ntHruX2k/CD7A2Op6/ZqzBW7EtOzPC/0fFEzMv5B3hOtfCzEx6Mm4t7P9eaQJVz
c/GFwogx03O8azje3D4Vt/XCGdeMhxNzMQ5SVYB+AiQinzLrnjLGXbHgeG+5ZH4wV9B2JbLUca/E
dM8+LcItXSk0tpKv7DeXMGqugo+4NwAKYNyrYmtHEok7d7jwLfcOtxwpeEyJnerbvUoahK4CsD23
Mu4t15q7blYrcGIUNIGwiAnuo/ktG5629FWdYQx2LUvpZMwaPbQ891qttzmEFL07OvSU8eCiHIgM
mFEKyh6UYYKyqLO/0XVRjRPw5tHLb0Ce/OYKO4b00rFdeiRUWt/mKgbQEz/a1Pnoq/ZmmlgdECz0
1aNq5cFAZb2gvFlXGDV9+Xb/URqjVZdQ3lQRtWrZCMk8izibe8AhABag6ozaGBD8OnV0AWs4Zin7
OLPYZxYYfeOmhpex94V/m534B051xV5b9b3IuU6WnO30kEGKWpOHu9mQ3mMpo0ReJ1lllQPRGNJs
bnQUT1o83S+/ZQzOtEAebbgUg2j/2WQ2K/JRT55P7LfpQQ8mElxQCKG0SPrn5AHiHcQHWIaxSSq8
JoOXrXQ6DnQt7lC1Go6cm/EmNnIgL/ohcYmfrIdTx9aM+AcAe0tGAR6FTzTspJS99JDGwv+QbDaK
l0QRATPIHDZCUCTJEhayHdpMGY1CYWo+3cnukvg9Of6l+z+hpb9xJjV6n2O21Fyv6/zX0pY4F/TD
w4m2Q28sFYOz+jlgu8tKteg/26Asyc2/dVSFA2VYWGJnPzbiPdbseUPmgCZkCUs3EXP1dMP/pKba
RUMefUMNUhHBn8Lu4JlRaeuneTdwBi+LtKmDSwOZTVNzi3GRRi3z3dUjsJpzMreOIiZ8oGZfIdtx
mVp+V+pLxYumePaP24eQD4o4rtVXUDtVM89Wj9v64eGJJvYNgoWcwTrD5K8y2Bp+bUL/fTzOxJF/
ehXZ/T5gAz1RQVPMEVCjx6lBXDVshfJGcq4Mq3TGT8Gj4BiLc+knmicHKid0sKaLCDE54FEswPEp
nCeNBSX0kJeWOHZNFyhPLoYlFsUNbqKeO7t/V77I47dRFxi3SnWlTD3x4z+88BthlV2zvT0TbLCT
u7bJPGxxs59/haKUlyTaOCDwuouGxsVF54mu2+ULfDC65nPcOgyROm3TUuRCfar7YTZw/yr+kcky
SylQw+LDHny+kbErtk4iuwfeOcq3JUX4X3QR20934V0U21Y56LS+5WtJ4e7ISk/cqGx395500KrK
Jgk/jZRn8mz3YiyxDukUEFlsiIcYUwUbxMirvjcc3KPDQMbAMyQypSacJ8gCo+pzKVNpkQpbRO5v
ccRTbmbuUUTlzNctIAKTSK5p0BiQ0KC0bNF7EfusFjwOZgFeap62TgVe9JgIVLPG01ofmF6eU7cc
mJJYMTTDWo6irvsm7WqLa2Cte+aTq6gmgkKrXQx/8yfIcijFRO4hAz8jRvxnW745g2GT9Ml3IuIz
OI5FJsJze6qo8ByZTu5li6F49mXcuwgOVZm30ahuePgdjZY00td+PEU/cZdZ9n6AuSuJdop3FlkH
AibxTOHQjMX/ZBDSxY4+F9QPZIHncxpXh72ujYCsfNb66pRTX5BRnp8EvBjOW7aGYnjezThK3w0/
N3f5YcGDps7KWeIfNs+wRWwut/6+9JaGobmhAKShQwDW5L1RfAN/I5oRK3NLEu17yz6bOU20/232
0LCfGTOs6KEoiIoqNOc088MmJwZ78qqRYWmrrOlfBLJGqQQDV2NnmNYOf72O4hOZ/3/CeWn+JyZF
ptQmz2ZCriJVOB84ptlkAbzlqBj9fogxm6RBUT5wJGGvDsbfErL6m80C85rDWwCFauaAJt5kIdMT
PNTwN7qiucRRljYcvwdi3tPts4Mrld2tOWt5TtLa3Ehzlvmgd35u8S8tm1mtJRc00qXgEy9Fn4iE
m/3XL7+nYbkXoMc/iil3S/8W8j/3R4buIF7alwIONmOLyNlGbkEq3wMxhKYP3oRya1kOGEIlIJo3
1399F+3mNr82hsDJA3EWFoVLvAhTBMFOHvbQUOAUL8OvD/C3vXEoWLZWpscx6LG2o0SEeLTSiZFN
La+stp5sF1UFl1IEimivMybR2g0wozXlphygnAw6/2Px8f55rklf1JndkH1iNuI3Yw5XqMTDTmgV
hJelmkfEVYe6D3ha1mi2GDpfvjZ5vzMV/k4DBc3LAfDScOylD1sLMW6Fovn4TTKncXx1eraEOVTm
fPPyFuss9c+vEGxXzvxsVExssCXWEPcaoGh6u+W9BWu9S5dGmniUmyvlxcApMyd3cOpWvJ3jca2S
u1TV9V+6bqXqyd8nXU2IuQ6dy7VXUmfXN3nOH/47WeVU7s+Lncfok5xwO1P5j7u82GssZLcBH8I8
JFnRsF0QFlvjzQUlklBAqZYoMZLl5ojhQKoiIpXO6xGs8BtYoYIok/W7hLk/IOd1J1QDTIe2B9Vo
bIBU/VHPXbvirnU+TVs/arPDSqB626Ea/2fvxEBy/kMAipW0r8BUqWch7PWD7nIVi8mx1WmiSlLU
jNaenBTQa4E/WuR44bvOoKrGEMIedgnkCDiLi/VqYUtszGOfUMfXY+Z+GM8XruhcK97EWj7HQjDh
M4HZxBeKcIX0GUwk/fO7wH92TdqdyzTC710ZhSrdjZMMY5uTgDiMRofyhHjfNh6ureItnc39rr0e
9RsyT5Z9r89Xo34EEwA9I1Vah2jlAqvAA17uzxy0E0FfRzwNFY0IkMB8FLkfLe9u/MWfa+V0pYCK
/6LmexHAFDeJP0wC+AYfhQEeuwSrDAdJHk0bJ1xUMLfBQbtnreevSoyr5LJeNa0L8TX8DKCEYF7l
+dAslGsxuvbwzKu6YmpaZB1pbkvpU6kJ5dFunoKwdUzQxoD+IRbmZoZMe2muXkVUvhacib7V/Ufn
yfsUIJtf6NRnGnmDn2Emmr9FLC0+TgQfA7hfjUGSETuVX+/21a5pBbjuy3D4QIpRhlkPOZmWMLoh
fNF/1JSj1GO+bWmYZ6v6pZpqfWd/IfPNquZcATbCA2rTCi3aP4AT8CxEQ0aTaF6/Ei1Fz6Y2kcNT
BH/0hstFOwLCUMUp81xoZmujAPpK/xWjG0isdAUcna0BQxXA7iV8JwvAjheg8LkntCmkTYmguEkd
pC+R8PIcVEy4B6dKvGpeZppZKsQilqcWV7hUtnZxGsiSE7dWvoAQ8J+1d3yyPTaU/7yWj6k4qLTG
sfVZWS0D3V2z5JFy708G7Y02bOFFakjthLTDw7wf4P2gbKcquKLUbAcoMvQZ1U0J94DMdoguiGDZ
t5OET9DvOFxw0Si6D/Qs4PHqlu3D5xTYeQUCea/tLasn19PyMbCJt7udjy9JbpIs2lVkepKs7lW/
ycTTa0E3SVHq3/53i82APMk3in2Gmo9XJO8YOd2WerEEOOqDiAhHsVzbbNiyHZWY5F9HZO3m3XmJ
Slx970Mq4VbuPfjl6kItwdpLVvWgJLUUji60pbtMhtzYuyzM+KF2cizxrjGmvpJBXuq3ryBjnIty
TuJTtVuspD1LwjRoSy39XBzrwauC5va0Ae7NBYnSV3VbGcpoaz8mZB6oL5iqf51kqWvfo2sRLbx1
0zBDz1xfaKNC5+mi9nhOxUsy/apYTRHNIJrfDJK4kqQaDxwu4eCD1MsCb8udHzCNE5LauVnu8yzM
C4jM7Zt5dMz6tqhMXFYI8qkw29kXod+6XpfsbNO8bSea/m+pY/4JxWO4iX73/MrQM7IfnMinxSfW
tmSTUlpMiH7Ku60oYMiwWCHzAFRXXi0h5xB83jFCRkaiRaMLMm6dZ9l89baV4z2BJIoNZXy3Se5Z
myXc+coAcVvxg9iaSWlXgmnUALie9hqDUGEVtQ258WPUcEXVR0o7DPoejSqiVfgvHbrLMkqsLAfT
wXwiQXn1Q7auvPRqv/IWh+cQqtd0EWArLlKtudM8QA0wL3m6FKysfHTE84QYPRko/HG4ej7sAd8Q
v3x5YtkZ2YQ8OlX7GOLvHMCYdmQ2juDtcwndlZFVVDLL9J3GLdaW7zBEAJf7rtYzsU+NjN2wzoCY
W2s/PxnnPZ/iDx0Hj1i9eErI6TtaxXnmxw4qdDqnBn7mUKs2tIhemCnU+OxQveASSzHEEmOmuArk
P+E0kVjdn0JwRC7SLq4D1jS41A6jSiV3+Csy1kWacnkKO3u+zd0w5YnuMc08NS398epG8WGFbCGf
7AedIgwR5T8dW887+pObM8qjR1r+fYhMsjgxS26BHexaxydRRZmPp1Az+Fo14K+Cz00dgkLr3j0z
oUiTAXnarxcmtM5G2vfumPYwuBG6j33rvh6CxTF7I32wudhBoXfjiJwd3qdaMMJ7eYiF7rnp64lO
21IKdXuIKp+ajqZYhydajUZWu2N52QU9Rf5ww8AzIoPZA2j+Ia/FBsKiUTIBhc77YHz+cC4GRYqm
7/fGxD1PNa7b1/fYOwx5tAMd46Vo/44sOhTpQL7L7xjy4JUuejm6aF5DvipoJ4E6RH88PLeUJoBt
aalHDq9yn22p8IkTXBKwzYLeA6gguTfovCQlS9DpimwTghQSR4iyD3OtzDqG2OPlGLbgSiF51sU/
kI30wPDJJIYk2fXLyN2ycXzDZEGIyAKF8AQ/i7iyQewQO6mHH8A80F4x3X4qihShf85EmV90VA1h
hYdDA4LyXCxvfi6AFMKI36PXXqjNLtbrd2Ks1xr8Fe/nJ0CRR+D047YZj038KP0KY6sPAyFgrP7/
TgkYysAig2QPx5N9ohZ8BiEUHfB9H9EkPKCGuwmEnig1hoHobvGn+NhVmVHv2hSb9Qe9+9IiNVmT
QuO6ePxSzwJWBIGO/9EpeWzmJLhWXtfp4etazuDccwi1slIzc2fwPfAjRoKbbCw5UynAnEMj75RK
rwgGAcymd2M/KQcp6v/zqMSK/qXkY2qTFTylPBPHk+FQbOLLLnEJWQ2/tauetL37JnxinXtpptPG
atqfXLA4NXZoViixYp0FnkcNyHCEBHXTUSdYCjysxGy4qhbwz4MbnZxF+5hukFlvLZP4lrqOuiAk
J1V5tgZMQckori2/aXjvgb7iVTxSfz5QAaprfE3HiUx1vjjB2NmEWbA7LRyJuW/dNAK1bn31iQh1
+KhamqOD/AV4mA/JXZfmlwWMDsbQWW4Q0b/xvLe8nb8oyO4Q07BLRntEIBzBmXijcA9RiG7Bgphi
73ZclmHLVMzCehh1v01A4H+0zPg505uiVAd1dJPvhU5SFRdRzabbJCyU0M/6hrDiDbIb/HyUwlRO
zZcsSngBlKyP41E0pjzUaJrs7tNLwYEc/JmqHk2EHuoge1ujJQRSW5g4aygJeS7WA+zcx12cd4Ul
BF+pMIm1ca4VxFsNTWQlIFNbOclaOrdipyE3V1b9BLe+erT5HNwxIDKw4Rg/iCGVfCfhAuz4oQ0J
j3VlVkVx6IvCSEZTeor6MW9z14lt7mVBSQDgenXCralPkqtStAV7o75ScVggqbCoAWiZ2K4f40Xe
kbJXiB+eoJY3v+m54w0fmPsLHRwsJWTGJsEbPuCx72mNGGhd+t7KSppGXfrYBlPlIeZJI4PcVEZw
QCaxr895oFoCyzfS22avpVOVwy1PAcxN6bMjq1nNlcbm2vk3+2HRXxJHcZsGgc86oBK96d5KtknG
lpoP6tSte2blU1JDOL7aCK6XkWDmmkBZNLGmh8V/w1pT/bQYNaTICnvLspLUFYKLifoRyIavK6jX
2OpiVeRgiYyZxspmexlN/ctmI3gs/zmRkvN05iwFstpiNb0nZO3chkws0NBzE9dcZJNNC3gU3BND
xzamkpJwLG7XH6D9kaxN96M2q+tBbxNDtqv3bmkGfZ0NYbyjj+5qz9gjLZFoovqJyqD59yKe4oeJ
Pl3+iCtS3TMByfcFH4HrwCRvR2YAtIN92OME5kveVHNE5RSZNZxywjMONJGIsKIV4PO+Z/Rr1cVI
6TT0jJee7ShODgl5NnXvunuznkRwYiqlTaXSfK5ye+zvgRTXfM1jdSnaWXZ8AxF2q0Zkh/c7sfRH
t44+2Dep9F9fwKqKQLDCnlq7orX2Es5ch3pKmKgpyXZ5X/TW7/m5WO3AziLhJ77BFxLA9E40mXQL
HvCesWRZkw9StjETRsXVRgYfXmUEsKEcXkLHzSsxFXOJAEV519vg0xHUR7yNC2busNlpB+Uasn5+
WdY8TmnJsHzVa97AWp+trVlJtJcMnWgjK7YZ3HSSGUEt8mIUq9XtsVnVP30t0K8QctoeGeTiwxvk
XlSJr8lExlj5SKfx9JTnZMl/wgzx1AZ3ATKgf+9uSORAWnKDEYCKk/fIABdIobrqSzXW6442misp
3skF4PT35/I41AC49UPZ+fdMb+LyilGAPD9PXTfhuCmkovFPIVh59mc73Ogw1EUaufZF27JAcjQw
Y/j/K6s8dxssmVu/1hpRw+qxsx6l/fJdLXIlZxJ6QX2yUWN4fiJHqtN6OJUSaGVHUlOsthlvVj3F
2MTVWn8feQAUjotYkQA00ScJBO8r3nW6GhEyJDs3qjQGTS/gA3+qkXKLUQmK9sZ00nSjZdRfikdX
yhKBkKsQbiU1fcSweFVd5YKBX7pM+Me8eSTrDDt0ouGclEsHwdXtluKpNLde8IeXN/UR/g6bl7iJ
03/Kg58VX2pdH3oukI7CXmbC3N8/6JhGMSyGkQ1yPD0yTw+hpqbyZZwz8yM+WVMdjdB3sG6FMVS6
gfyLZbJyP9pTH1voIoVNAHXYPzrjBL+c32DaxeqYhQCD4NREGAZ5QzbZ5f0Zp50h33E1tTfHhU1L
GAi1I+aSOb4hhy5NCzLX3KcKEmL1e5Gjx3h3Q/Z+Vx8wwtrA1PR6Tg8PpnKlGvJ0oWeFKTxmLUuY
MFGZ+3lmstYWw3Zx7bJGjW7nc1d7pB3aZ/260xsZ0HCAwZUEGXi+a6qsbte7tvM3swBgMMqtAPxX
hAEZx5x/U+Q48WgA/0T/Ztn0fIC+rducVwIm0MFkdXSlC0dbjFKEMVIkyiZkGReAy96zDpawwMVP
851Jgqao8/MlrrkBZ1OZAP6++HHzX28qgJ2sf9pbueWJzkBJd+F26PXr2ukbKCPLHd7Kl8X/lrrh
S7hF1Dtjx/6cfQ/1EHMPLypJ70jvgKRPkLxByv4W7jeBhyPjyANR2CxZE/z2OTdEpywP/8arjzd8
QxJyieK+o2m5oRsRUWI3Amf+O+uOK2GUmL+D5ei+Ze6t1KyDFAw8m3+vWHz6ZqV7S8lrfXC2NFU4
JrwMiZorI70GDZ9A7OuWBecGl8roqN/sysA00GL3AUzllCmTdvbQF+y64iTVO2yMCCWfIpes6qTR
K9TXEXa15tVMB+7/6pi8IbBxg0hh2/eAGNIk80cyyIItDbcxlC6sTF1XC+xjcmmoZ3kiUKApd07e
6/PfkvdPm0oNYKkn3TZiIkqvjGQIDhNYM+0k0nDKwR+cYSomyZqmzk9oxUjEDX1SwZCMTDlwZK3Z
bgY/16Bk7FsbCAocFIdFbVu/IuMSZanvF6rsAkBW50kxZ6Ze9aGbOzHnwVhvcXWRp5Eeae3H89s4
D3B0Rg4I48MAO0JN5UMgti4et6YyDKRmvZX8EwHiudAisdn8vA05EMaiXdQ7hs/Cylj1bH4fwRoc
xLFZedBMj9Y7yhEnWLDAYT8OyNOw/PoGQ3t/L1NE/moYIXs5yjUezgxA1LTCGK+fHU0AtloB+Y8v
/sgejFQMkCvwBsadWtqN7LFzF0qlAYSr1/c2Oe+hSaey8axTEh9Yph/3w46/YYL4e4yUo+ZSKkIj
iAhy4JeXxNViD/HNrrgt2jx02mrN8Bv7r5j24yUQIMDxf9gtm/f6u92swRJEA7K8ia3K14uck93e
p+bKTd9h1WogPAw2mPF69qQAYSxlf3hnlRRIQijj9rG5F27eql3zGsOFOZj6Q4SU0PKYm/eDqFTq
vM6MUTib0LMbkEXajWPsqcYjtfEH+CoRdAFblbwse0rrSZtANIlgIaeH5mMtmQpXW8y0w8RN6w7s
Ec4clJxXI7HyszEzpInBbcXlgwvny4+W25gwKBJ6zCjppK1xeWkVGAEGbuPUkVCMxNr8Q+JYuBW4
SHJAvR7gWnq2KB3R+Hiz+Fc7pYf7Vpi14W6K94pPPMN/2SvIPcesdZIDfYNusWLDEULOdKJy6wLl
G3AyGyPjXFJ+2WEg4vmXyAQdvjmmL7UjyLcRkLHdtynNliXwxLISbUTjEjreECbDzT+5KBiMsW16
HqJ00qApCVdUKPQ3HhmoxFVFM1/Yd9y4I9aXVrhf0i5IqWd9A4MDNNI79cPAsK4CnzeMdUMDDaxC
1SPZ3Gh/ncCdwCvkGgQ8DDg9G7LETkMh2kjcY6i0Yz/8uzavisOLOLtRjxHBP9YTycXHGaM3OtTG
7X2QalPKB6LPzYz74HJXuQSRzz3ks+32UPm2axbIfANaM4iLc0xq2oE3unUz5dYRhbkmj2cJyLv+
+gjIZwwv/Fa+kb1Jh/vyrb93Cv5So8Gqge57RT9aohnDDUL83l+qxb9Xp5Hav4IwtIqWX22deUJH
ZcrsnjkGYRMNF+UfPSeDk9zJpQ80nabDyFptjtq+IM3Gq4cGQ+hjeFdwvpPaXFminlVp+lqmgoye
UdIFQ7C9IupXTCZnC4C4vxaPsmrvV8pKpwGVFNOWQo8rB8WNCK7o96cDGO6+pfMl7/+bHiCxOJ21
JX9HtzIK+ZQ1yhdCqppfXXBMRifywHtNcwEgqoiouXrgm9GT6NrihaEKLGjaWTnLwpCq5fWciNIZ
bfBe7xn11fZGj8ikpAlzBtnAg9UPM+A1dknseslW5l5FNKnqWaYwP5PmbOlOF/xddDMdaU+rpuOn
/Y02HxGShZ/CalLSKiYgJqq2DshJv6gOaQ0+dXR3pulI7cHC+U+3HJCIGPZUDQZKenE8VseyZtc4
HErTPyb73ZnwT3Wxm6JfOCU4S/VCLmOi/9bJq7Y676hud7epcZ15xWHmShGWXxbKBX3rQtXTgami
LMdE5P497TdpohY01gA6j2siNIEWH+VywYaakLn6MFosWNa0sAk6L7hG5L1JN3fzYxCSF7Xm3pb3
NVWlTq4KFLxkaBH4dWaIevixeXebwmhKZmsNZbaRjaq6p+slkSKUttBaaqJhCkDegeautrJ6ZGOO
C3J0/0HsJQ030sF90wpjJT498yxwqAceidQ+oiU3U+qZiNprrsLmf8HfFWEg2FatOkaJSYAZFGgO
jKoLd7POAs+KOhUccb//WqjIgicR8FVkTxsKFrGOe/9L/rD4/KK2P2KmIp1blTJV2qiLsyU0Gl81
t1ymgKDqK/17AhEnACm01tSdwS37PpJJyDhdJX+1/pvJX2gnVoWZM/TO1Vn2oF19zGoxK/dkMpFh
9pVjlgDt2dQE6ICPzkasi+wRqBnjEYaZ/fywZQqhNIG1WucJEOr4O0VUJ5OoG6/ycgZ5afHSd8OW
tLFhvzwVZjtyipQYzhaKl7+RNGfoGTHUwIYccDP5NsFlQs9Q17IOcA7cfmSmYxiGPpGuKZtWvcra
QuObzmbTHMJZtH7Jz8S2CVjUKoSj1oj1HoIIVOuCHVgVLQ7RBfZhf4IKj1VJ3sPmAQyEMgKAIr6p
ns1UB2c76rKX8ORATZgdW+c235704iW9cLj1n+uvTFHXy6w8N+18mnhBunSHzfPDh1ybhjsyV2+f
COINrTNyxTypEPDp9Hlz68smVfquqBmJm5/GnVqg9SOil5NI1hc/th1QJJ9suNzd7Ux75hsc3VI4
it5HaLgRBq/OP50F8ivW96n73HH8QzblOyCCS6ehR7TcJn80yEMVuQuFy5laypE1kzPmdEaODUNs
Cn9tStezbAiQFODSujKk8fSOYQAmvzk5vKkM7nRXm/PLpDPFSDhuvvFhkNoh4naCFCGv1P8bCBP8
vZ0M5w0Uzg1ZjQMeRcUV/3MS1f9RpaGdFEvFm0QqmuQnj6/knC5U4g8lofNdPsrARKUxjk7S5wuO
hRmKuGl27+p/DYb4wmaG4Hr/vzcZptcJ0IR2QqS+ocqNWpL2i6Fs+409aUX+N+QdVi4b4YijiSDb
oheyuU25m0gAnu3sDIy8D8jhaiqYjhD+PFyzZ+Nc7QNgUyITF8eUD96pHZf7iSgbg9ujUFNzyvG5
mgSTyFJFVZ8M+3a6PtAMKDrmLyTyVs/L5VN7HYC0tCSu8p7u9nwNV2/1baGVl4Jc3rnFfVR1z08L
u2+JfgXd+Ef12KMM2jhQ5UilQ/FZKWscU85PzJ0esVYC4vhbq9yJIUWEzEkyD4os4eko5JTF4aDt
IMTAlq8o1dBYOfJHHK/h545SFqLCtAaIiLSk99fNIzmhFDXEEGcXcKdQxxH5P26hCRiFTvecm4zK
QOEzPEDjJxMp9BpQHWQR0MKYOl7F0U4GsjUnNBXS/gt4Rj8UTrScYSRKLW1tJ9fk0yFnzr7tcaMY
DnG7Qn44780I6RDBuZvUsBYCdvgWxLg2+vkzTcklJKVbYrDjPq0jsrWFGstZSNdWoNhCRlpc6BG7
18TtRvYBz6w8RkLA0pvq4RD//V/iaxIsAev60MWZx+JSv/2LGE7f+0KWYu3iW4yS8I9j73nIpwlR
HZbR6+u69A46qlf26lxHUyLkPrzHywHbGXIY6FhBramt+/SG09ffCqzB52x+yMwjRrqJR8CYUZc7
Z3kBxCZvBrmA2fzKiNFlsUPpcHjb6gadqgVqEMNyE5tpnd9cPiMQXusc5IRY6qzNDg/mZp0/6Vif
03E+EqqtJhCDlxnx/57gG62IaP+znT0UfU1pYuoI9eZNg1OjQ+QVcPztN5PyfzZjI85d3kX+nb5/
FioHBdYaFvzhw7vN9KzdDcAfaXoKynMIlT/Qioq5uSlOocVix+H63F+It6qeoPuGd1b3yNgkGcIH
BludxjRFsWtYuagIGVi9lcvb++89L8J3RNaS7KqiOdHQqn2Qrb91zm4mgMOwxGopR/b/08u0TLDq
66X9BIkkU0gj4wHdmdFeMKelBnBmJnp+tf3WdA0xa4pGUZ5hn7wvZeGdijkd7N3MIZbXX2u4mus8
k//kW8V3oNiGTtniZ8SiVwBbwJ7O/keltp8sevu/7nbKihtq2MjwArGxnIuLrX8tZTLSMlFiOyFj
Jkqu1LMwa2uHbm5kFcVFRlBV7dt47RjWHiaLzLZumdqKUpASlnWOUe8MtYoLAT0ZOPFCB+XfjMqW
MdsFPRjlGxHphAFqvIGw5yE8TFBKLJRiF19Kulh+CgonZu3UHV7eDNiiN8VVzz+xmX6o42c9yj9d
bevGIwhWrFHOq7C33z/+ziZmXSSRAke6tPrNdUCL7DcLRa2Qxagna6xTeFBuLHfBcc2q4C4B1CfK
nawIEAJlOefj3xytA+HXYmmayUQB2k68MOyUUrR3gY6MQwmsUcakDBKL4H7E9Cwzd4Tp217UBvQo
l8dEWkJe4e6/rD/NOGPC+miscIFzeCNdyoGkw+bi5isg7HbQpRFCyYa9mELLxvKB2Pw2eoOOp5sI
nBvIymN+T/CorJWcAD6bLNUo1Wt0ObgVgTc/GEYr9Iay14OQi3c5x1qr5oV+ymqmoUEHRdIxbkoX
0WMSvEYup3Aq6Ojd9EkfJ29UTBXxadqXCM4kdY7TjCjMF5mRYiRVZW9R9PIVo22bRS5XbcPuysol
cFCRYPDhfFnYU5BtSI7hCrlyPNWNane1uGSFhXSaokc5/gnCjHX7i/tOBgVJPTIkVmo1hIwN0uUV
A3qP8WQj0Y7AMLoyXw//r8Z0EDvztuKTDcyJCjM90OGRZRWqgEItXjmkZGRMlGFmo3sF38f/qJjH
yymESA+mQ4qMoHl3Q//GxlQcDqTfr+IFYx2zgwk1JAzCjBlOF4m/SzbhHeS9/ktou9+v4iTqAI1f
Dv48ckU6nNAsYi2uV4q9D1Pyv4rlTSNAxY6r7g/T2TAuthRWt+inah94W9ZMlRJoDmIG4DZd4czG
czp8QdZo4MZFHvHlFkXZxdXMaAQ7t+9ShhQBYz8kc6+UG0vfnqqprTl6KrES8zAkqyQcmHO69ysu
W0Lpt7hhBnJGAtZBSijVR7ayiBiL6GKYBgnrnjBTgj/h5yIDwE3EVnTq87ufLmoBH3HdRceMVXH8
uN38fGvyaALR7GBu2pC1mb0iHJ2b5Uh5KiRBJpoFm5OIe+DPl7cX6jteE54YmesBfLKnw+CJ3iin
ou9U3fFYvQCrnbq2w+5Ur4AAQnH670EMeV4pzu0uceyAK2DATz4s1l+taFpeG2WuPVDkxftTG7NZ
IQudOCOE/vZOC7FvIaymP7ZQMybWAY2NuJtcfTRS/n5rlf0dLJQ9NPczsFrHpLJQ+zuhCNADdYsu
9S9dEWT2gSzM+ZW3KMkxcL7lA0Ud41ezGTFXM9fDwJorQF9jTn1WTGBp8jRscl0W9EpSj4nPy2p1
ENDUVyfZUWiQKB5MfsuCcaBXaJrrdVMNSkiVQUt6rgdh12vu+rWm289aUXjnsSKkcG0t56J4Uou5
G/QtQSYg1ELTm24tULPsEtjAwS/zb2lyY7vc9YMz/pjobVTDhXlIExnSajPbrMPYigMbe68M1vgP
nQNgXMZ7oXxoQMLTf2mjm2oVGOOopv0Zrlb8J/0qzYq0jypkifN59tA0/GmtXYfIx8Emse0aO3Ft
+TRMYlBj9Uznd49UJZW8WiwYpyel7X+r++kYHCahH/QQJqANA+V5wc4HykdoSZfzgKGMiMBdPM2T
sTmC+T1xLUHC680RwMEKjSMWIV9Sdl89QadcUMvFNTDwTdSXcC7gPG1Y56yQ4m+wQ54HRjEcvyWc
YMysGH7Jcafvu6rTix7xgX10iCdJGiEsZlIdyNMRvYfxdUfHN5/0MZ8PRwLDjiCvUCZxvBl88xBU
K73uyNDjavNAEu0QM2ht4ZKpNUlVT1Gpdv9ze+8uPYad00oMog7MBOaL4fpafz42+RUVkPSb/Ssj
i+cqsCpQ8ryTVL+qvt2W5f8gxWBKejtWG5PQuaDcaTG+cIqplGB6lA4SNo9xIpbhLV6xk9+KNWuo
Kgjfi8Wh5I+PzRDWVKz/UHrnOeCY0gNTKA8ai/MGRJDaoy197dumcIK0DEDRjS3ouYF/EDMh4JaZ
98JLHp9WQBYj4r5fNeESwl56sRlhrRNYAx94NaTkQoS96gSMUr7M/VOnMzMO0kfbOLjWADgU1++c
nGX22ESlf3MOdm6oQPrdiPSAklHEef9sQx4GullmfTWoRymDERUotQFYcwcLlPzCzo4v/dOSa9Xp
F2pYSEsdD1fFa2i3vX8Emb6CtsDNQNXehc+Kn+Pt/PwPq/takLYOQgGJPl5CS3+nQjz+GeGHVV9L
BgHOrz4x4M0XdcpTydnA+PqUCOzyfs/8NV2CpjxJTkc21qrR7JqLKRSFoMMPjBrQ11/0fJ80miDd
pdE8uahg0Pxv9y4SP4dM9tuNy1xu5iWni6nq+fQh6ve1kso881QqwUpIK4HU2lRR+hj3lxMLpoP7
PIGbSa+FpFNwyy9GLlMgc32J59P/TRKCWwTIyBF1WkBxy7dzRyinhza5lM1c6LYAbSqNx9DZwtDF
oOrd5LIgYuO4lQqIZa6bcpPCWFnxx32jYIEXJHHOfBQV6kxtoTFrIRnn/bqq9oicu1KosdqKsAs4
bfoWP/W8KblAIgFZFzIqa91/yNdKqaGJPVoWI3CPaXs2R7xdPY4ae3sRTGBKUubmDnRWeWL5GoSn
lbD/M9x3e8vS13roD6CDg4IOM1ogDfbsvp6eTdwWhB8aYTrhG8GGeZD/8mGj0PT0ph30nAN7cg9L
8jawTJISDqjtVLfnqbxXq/rQuQkIxbg1Yd2gzA9Jar97gFG/opEsnn/uKw5wKtb1zoPGVG7OQIXj
UvAkIPp9ylStczR4KQl46VveS6gXIBgrZe0eGNH6SXu67MY0xDAkBfdkgNqsQ8mCPtUCfZH9UjIy
QrfyGG/5ajYUtk0w45h/1r5zOe7znzrQOY8BhBjzgbaxnFLryiPPBb0g+iFFEY9D12+KLKqcyz/R
k6kmfNNTZ5uqd5Wa94nDdflApkWHqcWN9gxK2DBNsG313xw/RAfBoVP63U22IjHXfH97u2DTYgVA
RbGnLhfZHNHdW+jaUI3wP3YkthCZRrsNuFVGix8xcvKptvWqL1MpMCLb16ohXe7poefzWLIoW6ZB
qQ9r1z0oktwRHVtNpaqwHBqyBEjPNL3fBqyoNUKtwfQfY3NxUpqVznhdJ9tKzhHLJcX6WhqF6Plj
yXcM51sA6/Q5Lpq+OuKPO1kfs95SpHAVZeRGCQkrxM2S/zaTqUiE77nuA+xIcx5LhuEudHs3zwiL
w10cx2ZM/odqCDqG4K/DHKhzObJT+vn634UnUHO8S+0ESu5YCjGIEK5WfvO7bv7rT8TiHU1tPkkE
/5KzUqs/AYLV5bx4Odu1o1jnkXdYXTn0xpb/KbjLFOba2hVF4peujz8p5RakfSA7kQ3kJcz5FBpn
p29PFiIahAs/7g43CLdtRwuF/5rOjnWbSKtjYKEFGxhbdcndwGwfOCPhQU5yOQsKVVRQouqhoDWP
tls1vwPoG1l8mLkyWJ4t2H8RGsFJdGnFqNcyI3yyEEHpMQJY3/GtLSjGAKg0UgQmQx/CWBFApH8w
So5H+IGVmSY8yReFw2tC5TxfniabE2mOMIG0FZWFLj32qTnd+zhWhyYHdBofrs8T7SQ1eYOHFm6m
cMvf0KDn1Ke5xDa/CPzoK74kF8N47bGytuYu2vMWYCTgIpNj2mn6NA2Lusz9d5pLUV9H8kdEQ4Vb
kUTkdSmXQT2WbG5du9tSWyA8xX+mIR5BX768ZSMkY8AWwwpTdqO5kmEAAMqmyz9+3I3pGCR6Rzlx
CCwt/wa7hnRs+S+5E4kywxw2KSpiJ+NpcPrXY2xWvHL+1bhAeQtf8BUGO7/q9Oe3kBK4pMeN8Gao
Hx08taDiiSuf8EYXeNATgOBeabiPp2p0tH6Nst8i9L3tEJliYidtuhADH96Q0oQM4sHsVF0eo/cB
HLQb78slIbZSoq710mMCVM0gHqnIJg+cRK9Lrv94gozqpPDmLGA5ewfW3PA2d/Qyt2NDahw2G64d
aCrXYqCXGHABoOt/+6c61bHNPvv+Z20ntLh00i6IyCCZK9+/7NpKA44CK5/2g4wTmAUUL1tiLxvJ
u+Dk6XxKNem0QuM3ZVwErFzgLk6s0M4LcBlJ/VPE7AM+v7xQeM+w96xBXjr7MftoF5itwZA+Dv9Z
BKmYE9w3VvyReu+BcDzimBUdo3/gfJpbpLpGSv7XbnuzSAlGSRjjvHbnf0sMQp/8Zdzn/Wy32z7H
D+P1dn9bgWCP5NVvxWgAzK05I6w4fEoqVxSIJN4v+TkqJ8xG8p17Pxhgt2u6mOABLOt5mbM4pzIB
B+x61jpYX8b1hnaHDrELcC8gf9yMzR3m7BI+5Kq3tSXzeu/9D1itgjDLutv4yyAGr/End1u/k9EC
FzXTtMxrgcjX4QhOprOi0m73NMkpp9DRR1MpJ2Ph1/CDp7PoU5RbptW2LpTLtuHHg6+2sSfA9AHV
j7oAdmqiXjpXdd6zEqIhpmWn1Kkmw07gjvZrpbC7CbO3uFu5xeFmZnDe1KEAq19ADIy7cS9YNMHk
uM7r+RVTqEsu3MPC6xM8nUQCFNIEUCdY4WaGiD+wxav/seC0hOqw69HM8Ah/Dgxh3VL22hFfJdqJ
QVJxtXH/UIighuRsYLzBEXS7ACNZ0K/9EuHkJesDCUd2O2YIs0h0q4lgvIxCPBKvEfyNqQnEPS+I
lcRx+PfOmdCiyKpKc6Wcv1WS3ZRNnFVly9mUIPifFwbaG1JE/7s1Z1tAjLdqTDvEAyDq3lm1TWfc
NCiluR+Y0BqFgM0+06SG3W0FRBD3kZRuO6Qim44cVPbZHGVq62nPcWpZqGqAVsHABquOUU9Mh9b9
X8z8z7eVsWrj1s2P/D8j9Ge7JTWYTa/OsB1aV6E8/MGzKqCyPKrHVw0+Xe7IdQNeeiIPzu0VV6Ry
r9pSrL2zKxxMu68F3mzrpl2Mwj1RWywLKbMb/ySLA/HeFsv7N1bqT3hZr2A4FOtdWtrij1J9r3rZ
z0htEAMiWujsU3OG6WHV9LI2T9ZtU2Z5gBfIDujXWlgDILnHkm8hlu9C6eJ7YWtSULhq+mIRSjjm
tX4u93I8mBJUjGCdjHRAR7HMBmSIoYf9VIhBdWOxi1K2btjW3tNWfvxWD3YxD5HMnmJO+tkjvVpp
mmtUPKqdiRvfrsn8crTrPygjleH42W81NBQyWOQo77cwB9B3V69aWXcTiwOi+KZlujFY+kcPAHG+
TdFNqfB2rR8nQgOiCkWih77cmN2hma1/vfxqEGcvgDSJbCKsJqs9lTUCHTz71sQp2niJnDlDeJVn
Pc3hYC2iHyvvQsh6ArZ2OECfd/fMXRN/MievMhxTpXcmzgQOeiDY36Qf9x8hvqMmq0ctHYtwvTeg
C182gGNSDFi/6Y2eLh3B/LrcuQ0wUaoNmSfRJwrXtYkSi9F5qPn8quIAFDAmxPwtJdc+/9ipp+50
DuUUUNYJtTWjCBQ32uLsqf+lzUKU40+e63etjZy2bqEXjxaqg3y8vvoU8SSytDce2JhXfVnBlfe/
+NU+8j71o2Ush0mgL8KHH1+lvyoNeUd6V/lGbrAVIbsfQjB2jjS/AJWLEEWUyPG5+x6S8XpMT8rb
kyc6wJiGDoV6Y2szjU4riE5un3MzeTmbyvj8fl9E/E/4EK0iJRePmD2YQr5qb0MS3pMa/g2zPsxa
ogkIL/n9euOeFJCLC/pLxzcCxBCGrpIBJV7amq6IDTDGLe5Mxq/qK3ZKKb/CXhjxhUstmhm3zvNB
e+YvZB50RYwzX/JZenF0ZrHimcSvGsy8y+NEXWJEQt5p0gRRvwl9C0ZOhj1/OYTEB8FwqjBqZ3uC
PN/oeOr45cI8XgZMOoTNSg9QpZPgzM7UgnSP6LTWrmX5QsdACEgaqyM85WwW3gtLikNwc2jAMjl1
Zu0v444sc2fXRZQF8yrt5MRa0RZIrEWkQdcx67VV1+RVHU4U5ub78uX95Q9SIe4Z4gsRCd2ltI0X
kU6Vy+w0Z6SOADNs8sCjk0g7w9RzQ06eHQDBEtBqxWrqtysgB7Tp8QV4RxbIaD1ZMgoVXN3tY2ps
NTG5tSaGu46NigyDsNtkMWRJfIKSqsgBL0B9smBM8zSk549aZscKUZqEz/C1URR4Ze6u0iqo+i2Q
Hbk8zoJyBXVqsumKyo0dP7rJfPP7mkoDTl/7x/7NTDJZzYII1MftVxVlkJ7Wq9nwLUO0ximCtPzI
+Q+UtsFjGmdx/o6XjB0maXHQC20RAbig6weiJZa+LgxX73mlKlnWSptob0qPX3GJjvTSklCqtdGz
RX1mZ7y0WkzVqIOI5021kZFsctlIR/2Ej37UH0rBjR5dlWD/cucgQF3SAGbuWmCuDrmN6fJyTxTd
PZQzR4X6xRMHd5neeW0eZMVrblldT2McWmvDzRsyYkNTFGnHnu9Z5cyvhGj358CZtnNKSd6LELMI
FBimxngLpswdsPTqgfau3zniGfIC8PHLTXi+yJQBP++WPT2tVAqAiYKNpHrkTsXG9YnqQ3EHfgc2
UrIGiSHrj5ETIGVps/XRpjTdbAxyNQErQ/SLkL6IoBC1JIAdWQFQDEKcqgnNucoZjjLvHa/a5b/8
94Fw5tY2FGo0xJBSGPJcjlJiPw6Ywm0AKKKiPBfnrQtGTr5IcTrohZfdaBzEgFcPfVu2TtB94219
ZI15qo7wWBceBTkM3eK9ders9rpmml1Zaf8q4EUm5eipoGPo7r0vvgOTz8iwhPY4KRX/stY4pfm9
zsJSElFPeEe6jeu93oXxC9B3JyS4jmz0VK7aA4gmzzCI645+ST3QPh/vL56dB08GGO0FBPuYMn7E
cWGeTNYWoP2mH33xcgLM+YDrfoTqY0zX49MSB06q48a2k6fx2QHtxV14BuQhEGtxZYPVS0KeNrHK
Up1/qYeSG1YAfzz7QcbnU6TZFPWDs3G2kIfUoRTbkEwe+1qEBOw00TOm91Tnf3NKr4JFsSV8uexH
yrQDHg7gCNMT4LC9/U3BbMsMT3S27IEY0BPRnDFeIHYYc6zUfuQvMbLLFys1QO6vZi3X9FCTFfab
QKHrD7jOaeinmzSP/0PXjx4IefwckwlHb5MYD55A6jk0rSHBjP/CnQmDX72LdjUpIuoUulw548SJ
WcwwzkW4SqxyYzEcFOxMuKExSkHbswZsV5VWCjbi+K3mAHMMTVjcw+Uk4Xg54XV3vxHZ9Jy01T6w
iUTwsEipRgB5eu6YaxzPQfp6AVRo0JBgWoPrpxStMGsDuHcbfMJsoxja5oJWhn8zncX3G7zHrr/F
r+jBuiHh+0ItXx7uhmWfCwWOmK7f6JEfgMnYyZz6kbR7a9tNCYexTe1LjARjNlpnJRSavoscFVot
5rxZsshW08KiLRDiPSdzT8jr1BH0vor0Bw1mPQGlOVaDCc5Gq+ofgIsBTtStVVxTAVnyAH/qEIii
IzBQLuss925VOIxMafcJW3+eAHJVA/JEpPIbQdqB+Ix3UeIXlwTF1+cGKtGPc4chJqRZzjuEHsxX
D7kE6cGt7WTHRFnThYRw+DvzETmJCJUX5SrMVNqObDT6a+Jc9dSbW+dWXNOudhXe8dyj1w8DxBCe
koG0vhbCXW1qebjkNYJ08DomSmq7VcWGEnFtLEdDc9jlCmn0XA3bn4+fgedLc5gs5NtH+ZySfF2G
/a0HXLd1DNWq+Ma6fb7F2gxf1yjRMr3CqBY3HlWJk0kNTJvWSFR0ei4pjO+s3K1bAbJ6HHJy6A6l
8YpQMoeEK5RaXrjYREDaPcNXrDabNdxhVQYM0otJG5sVSVYSwa6bhli2QcZ9hscU0ad9FQ5voq33
BQ9cIiHii74DfG+bWB+gki9osNnx1Jg2AEMSWgjWjqSgQICL1B//Cewh6iYKHVivY1KaF+wPm+a8
ZKJ7DBd18ykZg6MPtT2+F9Kd5HKjhI6TExOxkrN/xBtPwyhlbpWvzGKL1bfts4xPfZNguey/Mva/
59fEOpH1vHAIkNTeGwZ7HEiNdtyt9Qbjb+2kyxLlyqh5DmYQqZFxm/bzPTBNpdKv1iIrAOvC2lVL
YTRNWdLIW+3cHV4gJncEZNwCEpTB/nOOffDNB5GhOcxx+LnnJIQooxjwq8KAcecaoY3LYT4gDBNU
9yeR+UtsobMVvj7bf8PFsYvWRJQZPEVCrT6u7bKjqKE6OP3zV9rDWiQN5uPFCGmT70ebqU696HqQ
Jlnt/HZ0N0HMZAfOoIO0PnQAp7TZF1i7gy7LBI+6V7/aovc9T0rhXvZz46Hq0ULIOXikxoZhG1GA
thNTHkFpTozTaa3ur+ub34zRLzek4M3TF3S4G5yEz4jGcd2vF1C4r+QFPCypQOPcDjUvs+s0F5jj
1HIvhh1vTQOfQXc9LRNe/GPVER2vIjEnADvW2r7jma3STMs2v/34gbW3tLnSDE3SZQx9NamlQAlp
RN93efpG23j6ZtrnDVJN6hc8yrSm9YFvY3L6ECItlzl4g3VQ7r4FwPTOQrS2Sp7fChokLbbU0FJ5
1U2+cNAMHEFHRRrJvFIl7kY7W6FUaYUKl8wV9vb9LfMtsbWNhwCfxTAyW43ODQOaWIJxuRY6BuZS
cOQonxtLpSMBrQ0UgjUxLrPoUic4M7VGdvbq+gaTDmA/c74lOdZGtyeJqFhM9Kp4A9y6UTyXFgAd
EtPtjh5tPlLbkabOBv4V0IiJSiJ/inSl0KeHPnIvV6aqKll8PyGf9qEEjMu88e8iftW+OewP9KMB
At5lH/OzEookVlQd7PBwtgpPG4lVfcMXDXwT5Gj+wK+I8G65wRyozX7M6Y3+mzscV8GjktiXj/r1
nVlA8+bBchwx8TYmJeV91ZSRQp7M2cuHQLUY7jQxf2no2dXPuz3gh+Ehh7L885RhZ1LDO9L2/w6w
uZ+z8cP5/qvNc4frNEcS2E+wzIX6pbKlOxF0QrYo2rhB2Bi5F+zJAokXMgULGwlgbm6pZy6IXJgS
DBEzCXwjC8tszaD0ziHErm8lw4xMmlsR9NqovuaJbNYHJ64Ihuh34fvQ4+IV7lv6Dnt96X1BXup/
QNH+znU6xrDVDZF+jElRueKigu0ZGxGbETqG0JhukTr2VbX69BpdHY/leBvM01uVBypdZkDxdrjI
d9V2lshXIW09RP9Vjsi/gXNynMC3Jaknf92rk+RY241sir3iyqzQt1GqVONHlyi9VpCJuUtj1unz
ubiHfLDWHK4x7x2QUYdoe8LYpo8teHt9Q52yfy+gLqiHRyIO4G+TdI2ZqFMkNnekKShUkswG49sP
bmHIHYMOHNGxMc9h9H9no5hZrx3nc6erXppoOCFoZiqQtw/YXIDdr06BWQ3NU22/ZB7qRQD6cDmz
rCZ/kSPfeuSp5T1nBe13u4XEngQK+IdTZhSZwpSAq+Gnc0HxcINOx2N6ERtQXQKW62rr9BbeyWm9
cGXttTYrvQ8/xh0hTiMLxgV1klIgprSLkiIQIMFHyUW/ZsUemvGFTG85aKXya57VswQoEPUSYVsT
ZSST3Ct8vAEINonljyN9s07HyApxCBHL8cUVJ4luHeRRHVa/QRsNQuS8ACh2od2S9JLxGtbvKtU3
YLPV4jORDmi/EJXAxi/PdwUu3Mtq3WpJFuulopSPK06x2AUWwgMadZ11MxlDFhrCYa0F1HOJ1x2G
kPShkn7kk+f4upjc9IWcuL/N5JvhqwMedWwgzrDj1pZ0d0kVw0kKEn2yQRekHedfVbao/bsz2nFH
eV1lGgmQTX3GvqhDSbcTUbS6dJTdTRbQIMVyU8Nuom/iaiEoV78PaFUJW2VH/sMa8/lDEDg2Ogoq
kiXfBgbPwgM9U9oN8PR0tXtKUt9DKs2bRp7jKAZN1kBgPQ/zw6vTbI3IozSNLuG/LPsoDfNRvFGd
/nt8U1jvA6dzLuMS5gzmjpYIcOFIdKe0/9rpA6zoNsdmkaWC+wZh0rx7TbuSMNsFc1vMc1CIHSuc
YS5AGBOWt0WUTvQSjJQxqkMQWQZm8rhZ0BYAHw+6RZH3YB3/wAYTMdAR+WnssSF+Zq25l3QlLy5O
TpTJNk+objiKlVhFVBU6SJyct8931TZgB4+PkMrlcoC2vlOB9qko6TGfpVoJ0EXtcDO7ILm/Xj6h
4Ps6qQJt8AYnCpeWJAGbIKnuRb1pd0jDXXNykzDeqdTY/pk+Q/SwzTcjwz0AD9/tsc14xkxwvJQe
GvzuJECl7rq3lH1XFBiG03rYJTQPiJdCFff+7G3yrzY0TW1JS/jVUOQhvJVI45mmbrQl5S0v7wBv
xfWtg0a/p/WCWCZeRmYxVHBUkomsskklrhLehKOJR4Qz9Zrt+xzqM8ey8VwnwP7BvBe/Tvpk6W+p
gmG/flCeGqcwzG2Wwmk8e3zriMrpxTxLnYjauPHOqEY8eyFFZZ6ra3toT5xIU9MP7Ky/vCdrPuuy
1c9+SQkcyX0hxnc8lzKNcMpdcDiF4FOwQQH8NUBCzXN5fhLi21Zt0R4juDYjq1s1z1h5Z8Rm8+Mz
brVtsKlbrZgDEklgqUEGpK6Dy2iktNS1OQYqk2vOxPdfg0TAm7aC1LhAFS+X7F0Ai7Atx84KrtKb
PtncdSfIWA9yTCoqdITUgnFtT+nTQrWwe7gtVQ+gy4GtvuYK37o/usvaJ1tB5ngdyRn6xVF41Agf
yiP2auIGA7pSNtHbSLguX79TVFFcNFeiuPTJAuWrbvvVibYmsOzcU8OyT3U7sx/2iqNdSTpSbxP8
FimT/cTEvMEuHsT7ewED0JfMM1glzR3mSo2flcyaWtNu1uV3XO5rrfl9aWcdSldof8/eCX2NZWMf
T8fwM/cSqk7WfM5G67cD+6v36+rHaU07ldi2X6YEk/yhi10fsziOH9R29FWQ0HQimq5Et9j9fmlh
HnbSMCG7nMd6GJWE9Oqv4qSNC2oHqJLnp7jwZ9cZFYnE6Bgxc2ZYk7/YBs6fN/09YknyeDelh2Ts
9pMA5gbpYllxIEsIEH68j/y1cYNfIw36HwvFgeoO4m8CSkFnvf74WKyMqIlzj/PcilTvnNissmhg
gnRaawcrb0y/QQ9qCtf5ziKfKfd9GAzRy3EnL0rZMthVjtw2FwWFqOqJdXbqiksZkXJeUKTbUJyg
dMeDO/GBr3DkVEZtp/9ShjbnsT1H3nx5gRwsEQdGwZmSBxVeHlAt2AMYSngEHEZqwfWw5Rf6AaWY
djGoPigEn7LsVtNK/MJVAMf+1tdlMuacbTKIWlqKiBVcOK4KmYSMYI++b4CVQpMFy5jhX+Q5t90P
SnWpSLBX5wZYoW4fYoTr2sx2ayHDCNfyVypDBbdcNKDjFhS7gGFJzeOrzh528A89Yx9SYdsGc68o
YDedxoD1SdtINqLuJ3aU+wILj9pnSeVXyn4fcTnaazzySbZ9B/Af83YpgBguO0GOQUpOyd+9tQAi
hv9PP9tRbUzqXeM/KNR+fCxmH9+U+sU7B/NrLTixAEm3sRQoHka6DOMFwDBBqPa366NMxJ/xLiGG
bTmsKShs8ZV7kVPATV4744HZBfq4uiuqrjsB6Ou2WPY1jSehgBTL1uuxROKPgUBkLdtupM0bJrB5
UBXS6HOdZSbpYhHLuUaKZ06iX/rh+x9g/8dE2jzj6HlBFIxPhuT2JKgu97a1ZVebAGsrNXSK9sF4
J7SVflCIgbiNV0v9G3R5ZMYMcGTf2YkHCdXogVNCkBx35Q9SmtBscGyeV492xKb7eKzi267/V5/m
npW8NKR9Z51WVzbznONHvjf5BgSGks5mOnfWqcQfep2pTkEh1BiikgiuWIXL+Oh4Q6mmYH9f/oD1
MKVUF3wnKIOe4WZF3PmruY+/cM7B2j3jPpzY0sxDf0/x0gaINZ5j8kgcFZcfv6zn9NocLA4ITMih
vp7bbwidfQcHDC/3UzPR1elnZvKQQVW9qLVBK+XoYK38OTcxKsy4v07TNjPG1e3Ql1T3ArRVowQr
FKjbiViv/86uQxxc/HwbBBAN0VlAsCnkTF4q5ED09s5erAU0sOkpFnvtenCV1y4kFXRAZGDFZkwp
L43rQxyn4hTopnvB+XQ3BbDHp3ZsccSegA+7KeEFZrWED85E2eSGdnAQ7Cg8FweWIT6dMJ8CoF3V
paD53P91B5fntQZjhGjUqURTDt04R3d2zqIyY3o6gNokc/bEG03EhMPNATphF6IWtOxT1IgCo9mT
3qVnDAVkDVVOEbUdYTDwkxNoZYivTpCQWfDtBwd3a8R1JJiaVlPrFGRXvnhuFEMNoEq1BbPWoyY2
wKeh5VkrOJpo+7bIspxOoeJuqPnNMW6B8sCWThREyz3+MPc6Tgk7i9QF8gpl4ak3rpVKzLM5ZNqH
u2EKQAZEmwK3g54nUN6op4YT/zd3vrcSzzeYJn15C/l6HHVSCS8tr0Fc90jzkU8uCgzzNg1I1GUy
x1JTAfi62PVn4YkBrSOwOph+xpS+kjrfBQOHI/KHGjHA4t54dg072z6cxgH4q0Wya2tW92iqIGFU
1+L4XaoyghDU9WKzOwNWtJXIvStnWP+igZceFt+jN6RwyMWwjIu+HyfBi3+WDVj3Ekw4X8bvREc2
ABByp7+B+xnIIR10i09NKDNXDtkrsEBmIjaM/qMG6K2b+aQ4qgUOm1f3T8b21Fyly3rC+5lbsli0
jt9PdD91F5fYjBnVp1KHcxt1cehxLRP+u4K8kcFRYylyZNXn+B8Fw7JoG+rozRvoDMx2o9hzbceb
EeCZf7meJpIPfjFqG5K+rD59ahn39rDVfxIcZizHw/gzXLeTtAQw8C8q/HBVTDf+158VA0TTrrYZ
LPoyMviU+l4O80wL00GnVMQ6FOMBbnUuX366qNtEancVb5/kCjXX245iRiF5T99AQ7n7jyGcFQ8X
VPZXjoh48VZ7YcpXFAGnolrZqIfflK2voz65SPx4VoDTtyZYYvE95eCTiuJuTdkYuuixNvFMVAzL
HkAj3pf8eytVBabqNtClUl7suEVBvA9gu6nNxqlef47PdFwnAzFDdxzC/0Ky66vg7LarjcCbEJO+
ajBODEF8glJmvp6vsTdqV4nDF4LRukeFd4vCfhwJY9WzXBU26kQvxnZG9n8i8w01B+xESczGkEw9
NUMl+A+V3TFEdI+tiZi07p+flqspW+InXn+8xJVIHB7LM7NVRigUMFC/qHjLJKW3TVTSZN3SpiqC
UT24pFG98OGG7dH8n/XfYZ0+4OGZispWCubnF9ulZKVd9Upq00u39Y0ejDU8hOgWrdYhkFhfRmzB
c2a3JdfTpTWlJ6RxgH+Akf9RdgPc8mLeMZo0rQiIo8qQlpPFr8u+GWUzsD8HUm389eBMs/BE4NuH
pYq4vMZ6Zy/moesuWd8KBU4Kq71HdBb/uDhOse8EqIOzceuanfefc5T3j3TzPetLVZu8UHtdtKWY
US2tIxuvQrCZG5vXyQLj4cPTYgGV5Hpqd9NJMF4L8cB6uXLpQE7eDyCAANS+C+pEDMPrlXP5Hbza
TFbcs6oxC5VW0ULWELksXz+rgYQmcpDhMKqtS2it84YMAWwVStqy4ETcF6s2Et6Qeupf09XizZ6r
CWdWsAptNaaKNlkRJ7PciSMcDAMkqCnVU8UxsNgxCOt8u04ZyWU/13MCipwnIdBKtLa5uHwfrlVU
H6Yk0c6xy0+GSIUjSATP/8144sOMWKxpAw4E7jmGZEZEYQN8KmCO8iXQt+7BSe3W6BSDVwWw58I+
3CiDgNkk7aTvvCsVz9C7Vf4FLCvR+1BcGh636kQyotWjFJsIETGGQXTmZpd0W/KyzYLWoNU/J/pt
F15JCI0JHmKmtEhDX9T0UsylwZGfImA8UvS2C4beQYphhgSE0WB01cMEco3RRjM3AQnmErlLgnA9
ZK0epsdk63RYlesTutO8CcPixrAQNrYajW3B/cCSCvhipUE9aChtkupoW76bHTEiAHW5aZvliAgA
2qLHuQzyaOHCvWRdzTuvFiH6sQScLapfLiy7QpYoz8sc3vikPAvZF9E1zaKfJSALoxj4fMo1av/l
AxGRNBChsd1QBPpf7B9HP4fcz5ekdtOk2C7CABgXPDMPjiQVbkkJperczSHzQ1oLy31UdSME0tHZ
TCce5RhAjrraHq2LdETFjyydZxNXcZuJO5xBJwLC5MCxhgzvZNXc/oNR2AEBK1xSSpT0NP1vgKbX
SFzB/p+oUMci+rPG42ExN4WqYQDgsvSV/Ism+KDfCa4kOSlT/k8e9isYlR7RxKZKz50+4xcIcLt5
cIHQkK+0nnySQDOZxg9F7MOjDOU+NGoArDd8f3PCqeP3UPvzd7sASdESI9Ak4LmjyGKQWK1yZHra
nVG4qOPOPW5X7xHLCn6Ce2xRDn7v9KyNMdrzh0Gnyw698c1o8iFK7dNuFhm8zP8ZK5yU3vVJemj5
WChZtHX9GEou9TsMHKqkrtGn+NrcRp2M7Dn8Wr6ZhPuDE2oguWxuWAaoN8Z+PIkHJc+Xcwy3puRL
zmCj/Vc54DvxfwLeziRVBeiVY8RU/pfvs5HbnSDZoUjVIpz90itwdkjRRXIxVLqXle7Ha33h6zL4
XO+yBT4BAN7g8eBadSIDxWHh743ll5x1UjnYEi1e7qN/EuY5ADZo9EbXoC0kG8EfrvTxp+aJ1/xT
ee5BXMU2E+pQ41fIxJZduRl7gh0tFnaKplxXoUORitMiHqvS5voXQLQt1VaAcTE7MG72i+UoQFRa
mzeKLqOi6cBl6kLwS6JEdeblNCayezam4mwN3cM/y72Kv1ezPx0pe+8BNiHstosMdhx+R08hD8Xi
IhmA1NK7TO2jalK3upSSy4gmDq8W33rxIa8QuiaOU8FHbF650qO31yEenbddszIZFkyQWVmRvG/w
yblxX3GlgT0BLG88pasJrTFrooQRvXQovx5YihODGbDc5hIdx6e7j38CcnFuM2fDcPiR6y55HdG7
7QP2tQsNDfM6qKZz0jde4QuvImRh8GKPladsDdp2NdrSL6zEoQA9Nu1wmULztRtfqcxa3J4RZsjG
AxJIjCSb+x32W4c+VM/I0C8K1GArC4J6FcrBxEjaRnmFGeQ1+kmJn/mfm4xy+hEq/bddBWpFB/BK
+/ia68tX3GCm0Q2tDDp+SgbIUHhfBgbqLVPwT3Z7bpT+gGjdQ+d9S8PzYWDDMBKPIjEZm1DochvI
mHT+kQO9AHVe4MmHgSIL5r/J4OgtL0BtwcQmWvR+9eMeZ75P6sOLEopcOHLoWn6eEQnleR4PqiS8
PzqXf9i4pYvsWPOsVm8ZWs5SLnYRfS2HG6ZLLXkioXtbHHzs84liretdEKLvSUNQOBSar0MMLgNy
3DvHtcByaqrvyMzP1QWOfjAatjBc5OOYMSeohj9B8GDZn5/6WWRq7DMQgEv9UvX9VnvYX97YeI4B
zICBrALmU79r550d0lwq3X8VcKQYTGQ+EkFB9lbZJk6+zDyu9aIz0dKOcBKMbN4fvbhEeJdCPDgD
yC09U+TI5uo95wXWguWeSXCv7nzejz+5lfGWJDZ7h3JRSSe+C42Mf+xNGjvBlA/xhtgFMa2vvQYb
2lWuMsPwnwaHKkChqhUKHDRguGk77A6aTcEeY6FXHTioX1NVdfKZ6bEBzhb1Zd/yKG2IED5LUezs
95Fo0jLjWjH3mvYT/Lm6o+nMjvAlbau8eQpurFs7xDm36BtARNQswNwaO9griQdr7xAHAqBufz7j
PRK4xMjklWMKt5kJJoXXwxYL/bBOsShVOy1FoPw7gSMuu7JMOvmP94UZrrsBrAom/BsauFnAAaeb
W/5rJrW19rvga3k0eDyRfEMGXNlsN7egzvMgAWroMHq3Kg5SYH9JvJlVvQxfHekLm1k3dKviYS0W
dv3zGT6Dwpe1wGJ/dlKlDIujvnnNMwXDt4dZh4RXFIz9nlHcY91mQ67BW+pl5epOunkuXaeBMyOw
G4cHXeVYVdFy6f7hboVcbFtCj5avUwf4guBbkgEE4L+aFARDur1lMzYLR5vHPfD6EiFN3ZgWkU+n
cpE4wO3NbkVlt36mI0xSvQWByI3P0IhKhRLS6xNQKG/ZrGQhHjaIgdIlWYQq6gyhGBCqZMeSP0ML
oG0gtdLPpUpMv7KdneQUa14+VsJkQVZ2cE7NFrwleVaDqxm/wUxIc6qsPGVbhP0qfYekUJPXuEha
np8juTe2t6fuYiS0Ul6JQR2Jqv0JHvviORY7/idQ+iI+lFW2GM8p+GPDB1I6nH2fRP3739ijYMTI
nXLl5NUFZHqq4jqleVtP+IptHzAmelZKlxl/mQDLRI75mdOGVen1PwMBKs3Hst4EC5YhOtToM7XU
5TrM5q1q894rF2AKVLLAL659w4MEx9GuDCrNnH/FK0DYIhMlRwfjgqEKOO3YSUhPHsnbu4cL9gI+
5OyzZRH6yGu/HBYfDzhHVOaWvXWv5u1W8tSq2pylJUuT1fSPaJe2EPERk3QOSTbk3qmSBWD0AVes
GT/aj+3bl+1Le6wRla4VV1GUEpP7M9tYLfrsF4XoixLcIKsHJCPmZ38GrhHFk+Dl2jZLszeS2gf8
eQyY1bd2c2zlEhL8RvljVZ1cPWeYrimMh55lYjVbRsSiPepvfn8cR5dpFBrKY0VfccyNW+nf0X6p
j6RMTMV9NXf9FiL+jbtvQLcgpNCv7yMKRb7rmQkAEpmUyS37wlIivQUY+AkxsTOiiCfkUbH0ZPah
k05ZgWd1MZms91xgUbxrC980TX6kBwTW+z4XABzrlKQxkygyRXUG1fOZoCRsHhHyRP6qq7w4FjGg
jbhPjCpQS4biksZnfzGJbVjw9ZsB/pGfsrsYnfirGYLY+oOtXu1vi5MmNhsJWdlzvZR00+ANlypq
98MdESAZSQtqlsvDXsc9qC6HRrm7cU3k9l1E3ZZrQMRGbx9PNka4OmfntqAxXG3fZ4WEQTtL3v9G
LQiHZdA6gHcHy3CWcNRZtiZkgprz5370E4P+fb4p40E/W12ryf3+qTZrEy/z/bhq2Ci2ApVVzkiR
roa7KMiEwMHAXQCJhF/73lW2WTBBEixaHlWJ0O8kn131CaCXkKdLwNtlFoTootUd+jWa+/gbPXBP
xMGhtRUSQl+XRFqQ8PURtdkmpm8xI5ArAo7WfCvf71/FvSLOqtvDdyL2gewAQwcHgOyY2IY8MEyt
RG3U3IuViey8cGdTxiB7YJIzpGUXTYpBajgupPq6YcRnmL2HI5vRY6Kqe4FET6g1iJRVX6/qMsXU
8IYwdf+R7gifg6bPCJnwd1innPtBjVF8Uq0Lqht+h6uycxM5zTR8T9LqpJIXii0WdmUQxlfac/Ij
FEXPtsu4pCaFhXqTeRPVK0CKCOqVkNRbVKdZIx3/DuTAhaJB901O9LHj7JyguEgpivdbcjRaGc2l
zFSA8Jep1M6BphLn/S9ZMBvRX9ogQc4n8ulix3PvE9Y1tNcGGugq/Ipb92TXpOjYoJRcFAEHKevo
/c3gomQQ8VxYjJLGch2ALGTXJuD7unB3YB5ZUwnL03ywBNLBMndYUdCqvGVPeG8lhNks+dZiR/vU
JpkC2YRNis42BiaJRxfvyRWKI5UrwiPdgYtAGnMlT/s9lKf/PLBdOboC+Ncmkx+JCdGdbFd/NH1c
9svW6EjrXNtwka1NDUwStr9noM4isfddq8ZFaNl6RY5qyMuD6HY/IPiDdknj8hgXk0/Zp45EN/A0
gJzEBK1854S+GBSl6nQa3eqhTlh1g62yfXXSsixo+y4TGVWPjbQsuv04XOdkh+XPbwEBXI2HjAj3
nbP8Tq5/XODtipJvBScljBWSTXgRpWPUwONEtsZ81sNewB1lL369bbIULIAYku/9L0LT74gEq14Q
0xwhIUrLuewHaQZ968KLngDjBvyjcJxaiu8JFkMqzHKjFB5lM7IxREbdmRkmZPF/gyYN5BqxmJYV
PV5NF1Z9fRJwEwfEBMTZCg/3Tp4N1SX9uENGh/r2dlZFsMMiu8mau/cK0SX7G0OCqkAu40Ka+B5T
GalHEVw/yAYOSONN+3n4b5n/D6V1JAswq4DSRSptEuIdk4ojcb1+QweINFCnWO7521ibOKtY1wuo
fW5+r09raqTFMeOXUW6f3mTDVbjUbtImTvIKWXO3V3HV+tnGC2vUxPVnpIDzlIyFA5yooHgVGHRu
mPGLcTjG5j8K4h766gtSig3eUHDEfP+0/yOWu48wx1M1BqC8QqjLRAJLg+pM9J4dRSSHUw9ROTFP
eJP/dKvJUq9dNOun9R0NilrnDNMrDle9Ya320Tw0PQ9TEu1VupUizc2lqfW4qHtPCf2TQ+fA17KZ
cxJJmkJ+NHtRbokB9R/A1583kJufcGOQI9oKgcmOGEx4yCsHGHxpuYIIz0i+de80+CFG2efvOZzi
hNKcgYJnhOFrdHj2TBal4nHKzbfmk935LnYfcysQ33Ra+AQuyNxs1ONbWfsplIgC5RyQIYJD7Ag9
KiPtQ27LmAk0dYNqhkEaRmt8wwNr7bMF9/edDEbomCOTCoytw/byJT0Iw80p7cwZIZkLiEt1GlOH
E11M/HODeUDnb4i/kJVyg6PPcpSMIDCavTlVawrE1PPWiCMdWfsejPtnvMEjN8j/++Sp6Kq2p9qI
8ye2xCKYJm8jttEzWkP+qAHctCKfYIB7eK3ApWziiykg6fBa89zlmuUy3itnIr/GxghgpO0bvQVq
kIwQA8H0jcKr/FZw5jb/LMeeEg59ATeV4pl/fhZcleAfG0kXjq8lR3ypFogpd/EvsxHljmdwqUZK
d1ToQJwnwAXXXNneDHL4EnreHLpXF1noZfEz2QJANupY503HW+X5R9Spx+4rMyKzEM73kNuxfu05
IGxECJXrqV/D3bSZzNPtGeSmc4W53rCZv8M7M7e/QrpTn9l7MPmgUYnwdYAob5hj5dvYVGUKZdoO
B5rzi4sVx0QXMgHw9x0GKwGxCizyOg/bfgHM0K7YKehnblEtro+hMt7htkIOgE42SJQjAu4jBWLm
0n2PPxQB8QzLIKynzMV7Qo20OMLaGjM5OQZa7xqFotgbUpCrHjdOOqYRkVIgIn5A+4BhiLG4ZS22
rmifZlEOzty2MJ9XazwXBttRMX6lge6sS//q4sZKjeAwQfBGGxeoLB2kMp29mEMdFbp5hG0XnoYr
FtdjAJIc88/JzDkq3uIkrwk0MgNr4vhW1BOF7eJlCv7z0W8hih4CuhpLTk/RQEfc+tNmF/FQ1P9O
LWz/Y+UEeNn+dfHLxWrlP99vo93QPzeB6LO/qJ5WfyIfrWbN4Rg+K3FDEHY4M6Y96oZFiVxhQj/Z
gRyBNmAD49vd44iVeAQKlXetPY2gJxYVyW4vVfURvAyQJ2jhqSkWhb4Cnaw+B1J34lvVJVmO384F
lBmA6FBAa2h7/AsjU32cGig2yy1d9RgUEF/hezKdcCTUilRl/mo3o/zuEVcfPCyr9TxWAm23pvf3
M4teN8Kx962km6USZvI1PEzAY3Q60TbdxPfLFys3wj072oGhO5IVasolQgI9MGDxW2pCyTgJ//ed
xE/zJsOGiGDi2wQmnGjGJbVlLhIc7/xYNQrubXWdrxN46UttIyKJcpqLsCJWwGm3+vyitfzK8ZEj
X44S9eqZS//czp0+Q0G+nXvESrwgNoSSck+n3xnHvocAacAZpfLRaGR8GpTsSu3CoJt8UkriUdYF
DUX8VUgAY3lODb/bQp0OZ/V9xN3yNR34deb6gdbFUzjib8Ws/MXrGAsBvyqXj58PKnHRyecUDomJ
5v3MzfNejZPLLwlNnW0k+BzysqzXYx/7k5C8OL+oc4pMqMgnH3WymPDybvjDcbjsU+udpFCgtaL7
/RwoTrJ4bcrTJXx71VuPEu4iT4ando3wsnQIkQX/toxbOjVRPEuC4px3NV81sr9b/C8ABdUJp6SE
ojI47INASsSpo/OKfG+s4AcVp5GDwRSSjZ2Ngfo9O6nyFVYrHheYaH7p9dWyjl+oTAAvrvBsI2t4
iL0uz6Gw5Nhtf7q1YAE0ljMR7TO9HcgvcR/YGyJiTOZUyLdAyvOJt+yRq57OlOwTFXv6U4u+gRYj
bUcSBlFpEyq0DiFWCii6fsg18v5ttV3UO0Gh+G6HNk280fdFAYF6HpYC5SIcA58GtUmDJf0sG4PC
etyZAMyHiynWYZ082lJ06IttmS9rHd5fN7Q9fCXYdbaYaTJ5Tr1sLtSHe6H2hcKyAV6IyXuFseHP
UNydBe4SrHbLEiwu+/6z3+1JeTE5H4i75Mw7AW1jFmm7NVMrs2LsgwL0rj6yRWjuopd1b2tkKfx4
b3tp0+oJC+Z+lnUSYnyni/AtkDfypXqYWUNfyZMq2D80VScbdUats0Rmaw+CP6hd25mOcpEKMtOs
NzobXIFrnawuWZSA31p/MRDdvcs+opGH17Ic/DwcAgF3UTDK4H091ZpVWmQ8Rxk/9w+KeHlKxTwl
X1xblCgNLmFq9yfZvEQPewS7WKeeLRySgiWFK0ruHQt3AeEnmU9NOwj+OAXSJ9xf9Kz6DXUQdQZR
xaVRvk7GEnpyQuaFIkh7aQIJSCqhxgnCN7mP6fGnr5sLfOqNV6mAiwRKpsBLSrcj5Hkgg9SfyX6e
rj1Zl9g4sq/qOonDXZ22LjavD5qo3F/wQAsBndEnum4cj4VBwUGIWcw+8e4HJGAht+REyzln1dki
2OLPd5deWX7RlJ/zKazoAkua4gO8XHkWpMyiZ212iE0zH/xyyUDmgpNv8OtrIiDHIRdFGrKAOphb
cKnK82rnajFq3+U9FplDiV+lty0GLWioLqtjCIbOtOkmRQvE/HTkXkiNKRfiPPQ6P+i/Oa79z2Xs
74FjuF9oUtXXKMT8aViaIfHEeL6KEkNiBS1fU2llTz3ZMkhu/kc0rPpobdi/iFjUO21Y5JdMz45f
bHqnDjx6N3krtu/n1GFdvoytQUDG/19vjSBhf25Z5xNgATPuvbBPxn/rW0Zwyo3cGLivpWCZsgeR
jgO9IxLX8jmVgaW4eUMDKAsww3dXuxxIRKSQ0JBJyuk6FxOYaaJTonc3omI2osgFof67+9tdWeu7
1KpHwBqjgJMVHJlEEjv9lcfJDgGzEJ5oZhfoWQl5hlMD192GWkA7w628b+l4zjXv/9Yxb5QcTJCV
AS8Lb2OC3RF9XlDK9tOTPjtel2wIJ0Qosagl4tKyj/CLnAtFrrEb9UONmlqi09Eabrbk2AuMB1HN
1wZ+ZmAGwAJzUGht5Ol4cAB1dDqflxputR1SSt6BCDTYn6rf69v58Z/QSRg6MtZ1w8/HwIq9gprm
Tg6ujJzbfSGfeOv4cuBeopnib1xcXIyKvvao8Lwj5nll+copLtOYBVV4IsojLYImixM/rmXkjwRj
N9oVpeaEuwoEz9zI4HPqbo6u/hDg4Osfng34kLwytZe1xzhL5hi6rPVMs5sEpaPlGUdg7RYDsaRZ
WUXSiX7IwL/UqGb+f7stzMDqrbS2CN5/EoRhZ3Lcl5rzre+vFvp90+owYrmQGugsogb15Iy/Rznh
XnYNG8im15CRGbHTMZtXRP+ZtDpzN9iSqOMq93NGgpeOnNuwn8iS/wVsJjCQBp0yFrBuX1pyOHCb
GB6XVY4GLjliH1QDZSWw+CPuCj6tgf0b0fHh9O3zZPtrcwnWH01NE8v1Wo4U6T6OB+92yVBl1GFM
LFxkZ26a5hkOjmggKV7jhj+BwfCe3vqZ2rNrCnG4paQBiYXjhL+vbFRwr6A164srUqKCOYWQD2nX
wWVDsMUwV1hlkt/kPAqmh+0Qa29eGdpOZwvbJgLxVfGZb3wrfcDkRFMbGCTB1b/2AvGuRTPGUgUL
uGdqyrPx/RCx6wD0S9ROCBR1CnTW41BM8OjqXwlPfsM5G5IlDDEZck4FA7An0Dh4nNtVmPBJjsFr
xjFz16W3mQAoHl28eiG5Ux32olTEgqYXjxhLVsPI+RWD/FkxJ/0AqVGVFcTYLMhljElHpffDZ8vU
JzXo+SrhkLr3N+bNKpa/QkhFOhQmtASW6JXzMj7SIEZKxMQ1gUCqRqRh3hYwuBUVgVEe/N9wrlm/
2c1DINEGKSArP6ZjjsfGPhSFA7Zve1hY8VvIvdvRiZh+X+xlT5qGy9N2i99zXpD38wb82bHRfzgr
+d8zqHLh3yCmxd32xnjVLVqNZAB0/To6nDdro1DB1krCRH+wBqn6fFxy/zAaHA+254omgpApmt30
oXVoxh5hxPIt9MKNUmFAOmI2373kpUk9ivtBFSbOSRtt3CsCuGklnVO4eHITTXIGxYAo515Uw7pQ
1AJ9onqe6AHpeI7e6OVuEr3gqd4hg+P5ahaO1FZeupGNACzV9KfC2Uukm9zEx0q9ewIYMQ/ShjsA
OUQ03ub16qFEpT+Z9u3LZ7Qnkxs/UUx+ZMgac0imuWYessLAH7y2cJjvengT1sqHGOzuMMriYr4Z
1YoFoh4W3NQaVVBsD0cX/K374HgzAFoWVvPgqfk9j+Kn3csTT/WYeWVlEGLsix4agS96FwFcXxy9
jDlZjTWHKyTuOg9duyb7ajTUooyUsOc5iVrF4+NRqLJ6Cnc0MOkqSAxUYyZ9KhClhktQIJlfHUg2
ye8NLaSfSBunrbZIngj5dfwI8+80yq2UVov+ttPceu+b/E12NOTn2Lt1ScVKse1T/I/vK5YxsOEt
mCaMyBiHXUU6fcCCrGtHwzDZP2BhtLvfXCni/pgaQBdXsPVEKRel+nKNkbxcBVRMoABbKmskR9uv
z6YAGFNHhxsOZ5dQwBRMVuxOxVxU8R0n0OfKHR4UUiS/PTOjGCDKzd6yqYkzqnH0repiWTRgcaja
v2VtrX4WJUqDhG6eHlh+aupuN/DFTZqWAFi3Bbe+04JycyJfDQgDDXUUhO1IsJCLlzxlgs4NlTva
vT4zNpg2Asp775myVkqJioUjbDiAqxO4giPXpeTVYNehnW3L2CAePYKpYa3dEtz1kUJwSg1eRUhf
vv2lFfs97FMbE+0Q7AD4/XCRvLGroLR4Xv6pSRQmmFZcfQaAzFhPnBMosgTHnqywVylJTc8qL5a/
DLErgmFW8hFOKMwmy9sXfQKyENlAdM6jDe+y50Jimjmfbt3g2UnIt/5qw474QrPVhA7r9vQrZqVW
XwjIi+WXe2FltZG3TTyVcsqAmlEJkOAbPWl6fSbA5IWsjIw0PxsZW071U8IJcVhfEll3/ickNRWe
sSf3rzCZ+OX7majmTdA+BBplYpuRcRwjKASGZHqcmZMHgiejISi7CjhoJCLwZjQZzidD7PYBJ/lL
xxdAXF+sKgc6Ozhc8XvJAsUmOpQhPPlVCmLcsqbtVcHTqfBYQC9nNThjEUcrTrSyk4z9PD4G2arn
LPROVTQKr7NKYi3EdiFtVoQjPXKFdFWJEgLe75JKIN9Fre76ZwzwfyBI5iGRxSkKY+tXmTA6a5ur
JW/oQAvrbksquThJlaia1nzGm83zCk5U9S5sAELVn+FehdvaBeABQ47P142PHZHFX+WlouYyiIT3
MQslgSCCf9wCqRC81prPQfwlxtbYNPGAKXe77lhB74CPlz6MAsKQeV7fgnOlX9ieoG+LJsCgkabk
EtM4N26TORBMl+eQW6uxqdg+phklgHmLcGU/6vP+HwRXkenkPD0CJOPqaI9Q/qlcV5CkHXq/UQwf
UrwwYC7D3lRVieYFXyzrAbKtiFXl/FZJASgjNvwMNQQjl2AR0rgcJQU1fW/qPr1KEvzrqOEmCT8C
inApdiiT3PDxJzCiEn15BYdVMKoI9c195K+UA0Xr8jLNXxnCDviZbEZE4WuvKsLC811ERIHnwkUQ
h69zfawY8KWUB+N7xO5Y66N1P+r5RdcDk7e4BF4/NC7H49IZT5c98vipHCnHYv59hIWpss6VxWeX
moO+l4OoGwHkiZKPHJAJb1Jin16PYt5LPesJpwjQjNb7rMSNGbv9EPEehn7FYVzPawJ2SJW2vLYE
TyU+sQB+K8mr71ip95cMAK6ShHUw4SYiXv9GBGJlYdEiCcfY+CF2V2at7/uuTwOK9HDdExus3DEh
AKu54hulyvVIDWqHweFYnAoVOqUNW3W1UdDKpbTXsYJS3cJWcANfF4E4ed0NMxA1KIvOvDfn0TGq
Hpoaxstez4p5HNHmu1PSIb+oE5m1EQ5MYoiqw5s/0PoDs4ds9uAl2eBR29Gzoxp4sdIFxWHlS2Jg
sXpTWstvIWrluaDAke1otGCX2ghfnp5T+vF/x1myztHSnvoErCDJipEeIV56+C18jeHedBYHxnho
S71Lx1vx9gAHTqzAIjmX/iZGVL3CoG6EUbsGtuJW1zg03J1ohZ3qMIdMaAqrrO0Z5f5cnn8BVEdb
ngvck0iUftroHWtTTukTDP8ZwJcDSuMfHj7DdHotoK+FwSoBAsY7MceAIXeG1AZu+Kfb0N0z0CZj
o8CTMqp+t9MoG8DI4LltvI2TD3PkxbJKJ583Ul5qWb/5zbJLCCHSIR1vS5QiUGrc2wM1LUJj5kAl
WYdIOXS7wL8v8J/xbXvHpVmO1/T9/O7ROB03Dtm5CQUBIAvibKNQ8X113pCwB3lrj3s0a6rqT+Zr
tcDTC9xIHtP1Sm9reKksUWYCl4OHPl7+Q+K/WcqSgRn4QLKo4kNVZsmPKeGYgxzWhWjuHy4uQ/ho
mEniDLZ1EdecWHh23au1DD7RB34ERgmKW1Cz6YR3xmF2fYYZ4Xu1Tz2ohcilSZQxouOhmjOzla+D
MDCnN5E9RsjvkTOYaEO04AK66JwVA5zrTS/2z1zkl5PINEqWxnfx94DPONl5s49A2mTYkY3YJ3rb
+pKgvbPENJe5wc/xXcAmxJNTn4ukrw/IO7B9zHlJ+wCcH/HTO4A0OS5g9iL4mRrfLZE68pvAfJf8
FkzpzBgEYSXteeC79zjLo03Rph1s10zaPuRy52Pd03rGCa+ZQtZPKHB1DrN9316tJKCLLh2tBB9c
M3VMX9jchZmSjItqM6iF28l77uGOc8H7poGqHFpyyJ8W9HvTbnwRWFywZV+9pBBmscvj5i30uim7
9dgeH20s00bxf5TMEbRq51Xi6RrXdgOwQfoOxYceTneEv5O6/5em6MO0L6w6UWAYRu+xXlWbDOUE
Ol8Si3LZY3bzs0gej8vFEoa/mYP3JUlxxoHTny1UIuTNbFybnoGhZFAZwu8QpIEW3hYWxJ4lajpf
SIiMaL4guMRdB2Hsiq/MDZ2176zaj5exHgx/ULFsnrJCOHHGUXsrz9BoOhwZ+Vok033wf4dk+Itm
jCWNev0FTZf23WQJ9thLrTtFWFJYg7fFs5XuUiYS2BoEAhU34rVHtExQTtC0nbu0Izmf/q8AjX8k
QNpXMJitSGNwhjtWo/cQDZM/LaakZFqe4UVI+WkZCFeSxuG5rpL07Hp4hN9t1JAqZJe56ZguU5Yr
wUaFHDgIQhfyPeyTeXWgGjO+dXWjcw1g3xZIcNbPxgjcSJ03EKvOkiVW8vvBKPizhaq1kxJQLr4Y
FA37pfGL8v1k0ugmleumih8cOHfBkc3zO3hkMbYYMgWfehN2h253Jzf8H93LvDcexaJEfkfu9XQJ
9ogyd2H83zfEtL3hzg35pItH/HEkG1vbvbWuk2ncpUiPYGSYwjlHxoL5tH3J2a1aZjGbiEi/9UUc
ol6Tzask7b8fqNynGOL6BT26+NYPISRQzFdN9odWEq5Plgg8OESKr+mz4YSZXSnpe3NoUWHYg6Lt
QbusQnrk2vDTFa7lbwyEG52bu5sSo3IrNqNIFXkrm6RsLfMjTNp26X0vcIgjV7XVbqJJsoYb3Izy
dpTtpmghUJkpV0cHZaAWrupkJHJ0dX6tX3S41ORngxL/o/B/qthS+SCXWwYHtBM5WW+JMEfawbf5
7SJmMf4BSjHxpArkyhsAKMupgbBYc9VNkICy13vT21UAJ+Uhnlfm91dnage7Cu5cMjcZB3J0oAew
lLqszi4j8KgjrnbQvUj5zvTTWFoYnEwxK+Y84aqmyisoQAauUFo831nS697uDoJTUeocBoB0Oc8y
zfeo1INkPPGMmTcWmuPPw9Gd27+g+ZYOIBI8+GdNoRdR0eqQklejgvEQDkT31h4lqduPJ554AmCj
/9Wo7naF4cuZXUljZZjAp6+qApsHSz6hG1lrr+EFMOpAqnFjjrl9W9N/E5yc+gv3i/AqySMlGgV9
ISfuwT8b7GSrEvru/mVdw4NudRsvjDPEnXbwyvPwn3qhIuOWLiVPuOHAIR/NwLtzeD78RR8Iz5a+
DzPVIctiEEpCl5XWenDdnCuuAgnuAJQMa9M4q9GiclIsrel6vUMxlIUf76bRoQUnPxpBa8RX1A+F
sv9Dzdy7ZUOwnTdgx5PAX3m9PeXjjzzi8LVRkC8cT3T3m7ih0OD75TTQy8N0Er6FNhMDT3o6RIom
oeU2gXEkJCpZaRKMpArv+V2QA7vfuKwrvI99ZEjN3Ja3MeQ4gr7lB34HTfPd72PcwICfp6jCKNG+
asBNR91vkIwzNS6fLiw2ceSrURQ+p4srSb24EkycIezEn1U7P0AX09td+2w8WGZjIMcGXqrqP75k
I1+SL/bEakZug2r+JDkFPyESjYWlBeWB/+STpmsWhJneFoynrMOwsCP8v1x4jlrLJTJgteHA6riE
hg+ysS3UMEOSFonFkjU+NwMladbwn08qWPGKX8bIUXyvFsACoSyfKoVcmfg7qpZd9upUrk8KeqHl
jqcx2whcH0ZMvrk3hW5QFsXzm3mlFfx9yYuetKkoSkghmVntAK26Epn5SvDzzTY3Ga+Kum+y4+4f
52iU++iemEn6qC2YvsEQUkX39pFly0rDckl9Kuwfn4VwdT1dJeuqD1fMSVI7cER1y0AMuYSbi/Uz
JMPadtKYjIcCDs437zsIHzO2prgEqKlyBwkTXEdDAtFMLvBRY3686vhaA0shMVSf3cch1M89nCKY
wSxUjl8Wox1EdGvXap4uqqC5RFlXr6PEEpO/cDJbJpd6yjfSKfbkeih/Dl94tzy2BSWjsyxoyF3+
TbgVxeFnq9A5J7hPZ2LPSzRshRBQtxbFh3+GduoZ70OWMu0w4JnAaxse0HfBw4zWkdAA76hkE4ci
i23nIPypxAb0lHd3J6bu4EFePpWKX7do9ZbCV9RlXW7Uzm0xcah2/9rmV0KBYyvJwP+9Ji5W5zNa
Scw9cQpLR0raaa12HE3itjJnlFcMbCYlUD1pSFoe/fgaPOAtemqBV/2K7JwzlyhmEDagcq/u4Oeq
mNn0aZZiTEpn1Wjj5xExgPt6N6xyb8CdUoCkrPXFoN6hWcl6G0dHlWJ0z+CQyx3PYZFUtXW9Q2CG
nZdBxZd/9vpNAZELETgF67uPL185mUdikY5Nc7rz1j+yFv43iMycrGdtK5/MST47aQ9+M5cBj0S2
F37BBc2Qan42tY3lkKlnSgON+RN+mds8RJSaOJLGpmuhvW9NiGcQvNE2BzDRxJzRY8X1rar/OJtu
JPXclxTano2NTPE2lU3JZ2+Egpw6BUeOPcvjJH39hq9FS06qgtekLXBOSUn9N4ZcSvAHtXtmzkqe
d+2NihV/la2njioRdnadDcx7aNqykWXtMb7xNdBuUSKujjc1Y1cYdwdFgtA3xZ8CuxmTDgeZw9gT
XOpWH/AxE/WJ9vDJoaFyIo4tpAW78w8nGuZKx3Lg9IzY2uevMoh70QqS87QUiYIVeG30J7tfkQH3
7A+tP+vk8tiyd81fTk9lJQpZBA2G4hZB64J6hG3tqVOgZa7GTiGMf0+2vglykMRPDKVspoBYnDhz
5iVhkBWGQBVeuxnFjBq62I53twwzovVgMD88ezj7KUqW9+Fvn0v1hzAt8mjxwCdGHLUAv2iz7XYF
O6hrGng/Y+EMj6S9bOuGObkYnXYHR6cng2v9VLyefOz+NMRP+6IASGEpU6KyHDUykKgtp/3/ti69
SnwC6l0bnN1U/uO1qX8n3mOOg9AirasnGEGOOgNfcjlyzxXaM4gKgXinkVU4WSxecVIfHplDHwH8
36ZkhrK7rF9P/jg3rD/cGhBgzJ3IwbbLwYbB1TYw8tbIOrBZVEGyw7C3OZ+iN7wlbaWpp0StGnKY
H2fQBVy8r7s83Jw/BGsZspzLTAUm7s4cKekpE9Vbc01WhH2WF4mpMLIHrMWc4ybQMTUcZYpAtq4d
9tU2Q5tRE/ulM8mm4gTuqG0hnPCAj9JE5enNIUI6VRKovnMyOQb4Ndhzfd1/ANlbv0uveBloQT2/
r9yo0t1/ChczB0TPW6u4fcN4flEq2QsWxqd2xpA16Q4jvS1+l2LiNdSglNDJhveaKGK7hmrlrbEL
+rmmwdhqqZB6IVhVAHjXLA2DAN/AgHm2ToQuoSwjzi1XJVHL34VI4/8c/TY8hgbMsWtzkja9AFjw
bky6CDZ7F8lsPgvz5gql8S+e2eJHTeWx1MX6iAhjXaoB20n72tkrhaq6dCu3Anrn1OXRIYlcnSjA
CKQRDepO4onl5HhOWslxFmVaP6lp0usU0/eJo5rKoundR0TNDHsUOEfNGER/EM/F4vDpFNTXoU00
D+mzoqUQsap+O5uBVAQuUMAScG4bP6JSPhPljsZilibGu1+cvKHEneWTQTCds4zCZMbZXw3vxlhQ
ocpY7Evj8fBYb+PDeB2Pk7LhcBZ9RmpNPqy0cuap0rPkNdM8v68pERQuqQ7sLd/ZBr2S24XAstzx
7WPI7ShpUeY3/n6vH+P+Sd6CrzbjeUkj/5JqvY/tN2GwJK3ub4hPZA3FNQsu4z2/lXIlUMIeRhEY
p4ZG/PK3u6q4fhcsDcpC2eKTOUJNZ2VMkCSpYolUi6yj9GVaC/15sqTk5MY0y20c8Cy8mfzET7Vo
kBM0lXStwKK/i8Bv+nIrEphmXpzLAEwR5cW7iJTZPI6PKHH/qaWYk8Y+d4DfGCw2+smP0KQAKEb5
v9NWzZ4fAqzCkGKe+iGgHfIJUc/3M8VbzJK/JWTrjqLZP/KQf9c/hPn6Zzi+WFi4c5KdoZHsBE8f
ghN2N6Tq85nRHkZlz8fC9UVrbml8IYa1laUnRDRcfOrfN6QqwHLR4LUifPCAirgZ2yD1Gk2jPup6
Fmgy4x2hEovFltflyFBnAF4Y6le9PRi+iSOHOeF7Md0o9Xkuqi2E5aUx0Whn7125LdZm7N3tZe2X
1JKGxxAReQY7hnz5fbLDAUvLgJQl91/0k9kwca7EhTOEMb6mluS6Ewv5PDN1j8gS3AocHYqfPtj9
IQdi5IvEk1HNvrGAbaGRikpobFXnnMdi0/XQ3FeeBdal3cJyp7v9dtIH5iYLJ4YVWzX8Uj/aZu/F
ncewAaZzrN6WX7/Ilb6Xx2HEU+NgcPgyH7cNzFvA8rsNLNM3+cZFzyxNq07g2w/rGg8O2sKD07Dl
9CS4jNcHMcquULLqg8Hnr/3HuT2rV/ROmfhYjz/IdMXNWilq8OsG3y/NVZMHlx+cXG8k3WMlKbSs
RbqJXnZ1+bmbsDWuVQnZxj4xIoKpVa7L6hHvzj2MCLKiPm8RQKN0tKSIo4LCOulGpr0iFhFeu3xs
AUSB2rNWdAs7nntB7rN3P50y/tgkmK7tlcdxAchSkA1YM6pk9Ni0cBWZj7AmQCJiwYQO1Fv8+Ubc
qg84Bpuw0OQeg6ur49ux62b4FqPn7Q8+nmnBbiafOk0+E0nhYvPjI28SqAgKA4n7xJkQTXiVk2XQ
pMmghoAOXOfsnR14bf6HWjBz/HOvfGVW1CR5+ze049atG/wbD5xGWiGgvmmZSyQ5XQnNFx9RLq/8
WLY/XlZD2FajGnUiyCv02RdQqXkj+6OAcypVsGwE12iQAAq9xC4ul/xe6ue3fTk3HMmxN7E+8abH
iCysRC/HA8FJDdrJsSJOI6prZxe16pzuJOuD2+brPvVL34Q21ihtWQY08/KpJ/sXbgR5Y/vPSopi
HAOKSA1R8hXltjUNiA2DL+Wybh9E7ZWaDI2HrBZUL0tUxiSD3Ou6PQq0IwyWWmo7JT85kcsxu8W2
Asy/eBK0soP2XYdOyugq6p0a2lwLPFuw1kQ5zmshWcpdNb3rXoll7N2FasGvXEXyEkziQw1WeHRR
EuzfJkFfH+i4TLyZl9vEKRlLQzc8XX4GebVN5AfwVjwAdJ4kq3XU45bPOOK6mVi/OykwJgQ9wayK
KVLurcNWkPr4GMnQPsPWWtOrp0o/uqWrjQzyGJuB9nE1PFguRtN5Ma3HrqFCLFWnOX/tDmVBn0KD
h7gGAkKVNn+rMMg0vTzwZUoH7A9s0lBuDdTx/ejFTO2X4YofIfsrtLpZiYXyFpFp5IhzH3gMDMPB
nyIGqiwZmTsFb0qq3cLRBSl5hWqOMiGYkto6jCfB0FHRqWAYQvDkTSp/w5iyrI3zfGvMCqedfVA2
h6ZRdjoWB0VP/6F93NrFBuBu9PkqDqRDJiNxec+olqfhWTzGxNcnKf5g02F74jlDz01Xoww3E5A5
kh5v3miN8Ko1kwJUJKAcUIXWIWKn269sTp/IPRitypwM/JoIrz6yWI0EHUEBkbBRUNPJ6aIvAHwX
KF8tguDCkF4hQ8gjFiA7DRfkrKnbtoMShyLCW9RZt4JZD59BsDXi5bwsfoT3dq5nkABfQIWPnI7n
4gd8eXyUetneEVsvg5WrQ3SHrVq/rIUspN9MLU2eedZsQJk9A1Z3IMPuIOLYsOcPbDBJGSfj0Efb
0IG6SjgvZE3eH1NLI6KCHWhf69lNZEXCcWLH8ERv9R9RyZyHPtEMpXFQpEbGLbjJl/oTCkJHabyu
DBMQECI3TsnH+C+Qcqy9y0UEWlxYMhTDjC9Y0zz0wk307xAoSx90Nq1iLwCYcsydpcFNB6fKwdZc
qbA9neWQHNhwxRJZflNzxniRtcD8tZsPOf+IA6/cZBUDIBGgCVrakkRM+pqTLeNU1QVOSqWgoKAi
hE9oWFxbkWXx5vVrtEoCBDfpd1Ya/2rZjsWTkD8G+V/Z1oXWAzFMjhSCyaHno7mh8aBPx8xVN8or
jMHYda2mJ+08UUYGJXWG44Mx1FdZZ2tMNIka+Q8L/eI16l1O2y0UP5JoK5Izi2Q5BEYO96LD+3J6
GbunDeVV2tEofEPsS7cxy9GIH+zxf1Qslu9ZAggdV+55aIR7SJZ92Hgp+yqrj2SB49mt2CWYihux
If9chBppw7cgnScowIjA3m2fWofeG9IFzr2PqsH8MuYnbs6XVDBngAFEEV+7LRxjFX4zoCQGml+8
jMEbvY5Bso/DMq/wVZMKFX9Rq+cN6a2Jrw7LI8ASydsvJikxKKHOzrrn4HtvnvfeJgM9xivocoYD
hVb6JsJuY3iwyitWY9dvd1E2Dq6/NXYsY+sSmwnnpC2TRj24LrGP/1BI62qTMBRZKLozkwXYvHDp
OsHhFaC6SEGVuvpSqOf8OMLZd/4xvGJdsaITR97HlzTEKWT7YaBCu7QBRYa3xGLSM/VuhMp+6KAK
JB6umxZKiVu8BHWj0I3mNl16bo1CymmhJrifFvIpJRgaDdWEEETjh+e6/wn1jnpxvYeOGh3eZm3m
OcOHq+dk/SDHip2zmDF2NN0fpi0oH8rtGE6Oj3xrk4ueRE6qf9MsvD6zsdTLIA80ddYsE39CAID2
zveAGCyNu8uHL+Ek4JtxNreoQ6s7CnQ98dqYVchuciI0R6sedm1/HhUmxon25dT542vldKxHwazB
gwUpfON0MTxeso2Ted+PIfVfEFNIbq7gGYzM+S2IE/M9D5G+Z9+4yfN9leHj9Jaf/itWV9df8qT0
L3q+fHYduCM422zFYQeVE9RW2LrnSlBMhlWa7YCmLR69+pBgr+CSpfG8ph7yq246Ku1OTJBdQGSr
am5abT2xTEjBpATPT/0RRgYzb25al7XRCtSRldLkch5q7ZlH88WpE6AM4z/q0k4pVhAW4VBeXrSq
gnNgxKQKH+vS+HTqoRKZdpbk6R/0iBfRuArWgR71xcv0uZA8tbXmvgqheF+v74l4lRbjV0jHTR++
9IdmmNZ0aLsW5WH7C2luPJx+P+2KU3IAQjnfzf7tV4ac53qASiYBZp9xgEAFhHQaXhJwCosu+Gqu
4hIkP4PNfRPmca4DYUDsO9O4CmpLx5akOFiEHhuNBIhBMmXaOwnPVC/UGSJXL0qyUw1z2PKEgO5l
zcPpxNHhIqt2brhZ+iGzmQQNW0Wob93CtvKrbIUovf2U/0cExrfIGXrvxc8zx4hgyFIJmVmsje7y
KmDgTeA98IZPGt1KZCUdxBSnMAv/tb3Q7hKQGeAj+4j4yfyOH0tpfTp8T8ke7+fz+wXDBlhKaGsh
pzVCij5JxZYNitSgadPULjJuadUAXZpm3dvimUoPSgCi3e5VV5zNnDuEYCXoiCUqP/UFdtIOVyBg
bIW/BULVRKZpBtXV/2qpfjTLjTQfZaY3J5tI+CSTZt1xutgUNY4EQd2sg+CuISC6FooB9KcJ9axK
BSAHdq+7pf3xloPVvLT460INWGAgKZMGwrkf6nvqNuMd/VX+fCLS7Jy4aB6pndCbl/nvpaVxOCmU
5bB23e9Vx1NgCmRWXHRIFpE2LP+a2QguKhnxQMBX5jvJLQT35fgLxT2G2uupRuei2wTH5KJNxI9p
uE03GJjQKnzCDdbatki3QQ48O5l25qh4oiyazYduiywfBAhgL2CjkovzXCh5eTq/f7TlC0+Uy5Jg
ABan30NVxBcBfsrbFUklt1wgJrLc2EQGhgKOl1lX7mE9g2hx3JfJ826RfomChDS+KWYV6yBfNiQ6
IxC65G8v6UYIHlqDWqWzDk6Tf1G4/zFm17+H0zkh40utj+tRSSVa8cdrLBVd3wuFD+snofSCMrNW
nvQEHZ6uW2wg9Ez15Vge0Kz60WzjNlx0iZm7zYRE4FmNGRAX5yiyCWgf0dph7LkUukdy5Sb3kZYc
+6QkvDZt5VcQ1WQVXFQooHQ2EumqObKom0WL6Xl8mxI72xcmPrTzM+y3AO7RHUbLx2Niw8Vi8ABM
ekOodKAGoJ0fo7iSKf+3a5kSQwb9ursePp0XIZ99ALuxZJRYvY9+UylHLYIuKkC6vMwFisXGv7ZI
XGCvWCUZm/oCVo98kzsVwlQvQXGi4aRzWSfhw1iVlAtUyL5/z1as6xjvui8N1tR0Ux46xB4DVKH8
ss3lqtABAMTsuZKkCoXsmKdBxNFjogQSWyVU5/UGe4dncDnG96qwvcMHqO6OGeWWP+bKP5t/iyfp
A5Z5VDnirs7hlQV2tVQ1CBd0jAm7upLkrQJ/UF3x1QDIx2CrE2Cb9KnQ5GrGC75Lj7qruRxWzjV7
NVv48iPRWAZ4c2bdaHOkknlzjoIqs9pUqGk2L6HjlfrLYUPaqUrl5y4cLrC1JgfSUt/JXk8vZTrz
k0z03LNZoEkZBiz8lBljJPojqU12dQCFzYX82Xnoc+dzkYiKGetwJLOPShVRtKyQPcD/Tn15rVCJ
3FNlmgrTy8+5Y9mMqukjoZdT62AbDbhIoWzv7GVpWw49Eh0tHLVWXby0T9JLyhphMWHjC1V1rTcI
G0oC2SordGqMUy0eiD8ey8WE2kXC1Io+df6MGctIP5mgvZWrCsQis563vZUmZBwhGXF1ygf87GYE
9KogK+J3ovv7K23ErWldoXt/xs/3jSPe1GMEH858BqEtTa5ujhf/lgPP2ZD6H0Q0pmupHPLGkVBr
BKjwDlrCjpQlmjmvK3xpfUInnZwRxaAr7MteixDQgSV3OJ0z0hisplfXkFez8IcOClUJyL8WK9h3
vHeRLR2jixTUzdJ7r11ikPEZRKKaJIm3/gBHLeykGlltGEHIBP32f8h/Av3E8/cbrr+1LdxYjNqj
Rfr9i9RagMve3d1WunMWKScXkP6GXRcRZLt/Pkfjes+nKuB8Xmg4BBCM5+pNcuLCebIey4AOwzFV
00HsxFCjIXmyR8BgrCnhDSmr0J1JLZZN0qTzuXf4fvuLbe1WTm9hCTQczc82atG0NyP4xa2tqGKa
1dueecw/fm+BSlpgdQbeggyDNBIIIRcbpZOy38nx2Vda1VTAYCgjNXlzEVU/jrc/TG2dPsUg2ua/
ij//PqFSEV5T6/sxXmsZNwX09RBhZV+TKSNX2CUzamBqz1szfBads5vqSzbSU0K18aDhP4+n2Z0s
rWSzWroej7Wypdcjlo3QoWnNtsWd4jxO8aEM/qV0attZO2dTXEg2WXBZYzorzn1mjHqo0cephY3J
88pCCCzKyOgyluCmw3BvIEzVLt+FC6JQhUKlrPZ6jl/yAtls3hsac4P3qlZm6Uf4J+E4c1t9wOo6
9DO3M3H3utg8MtNzsat4jCvYHMq/M9yzKmQgyhtENShy4PLU0aaF/4Z8PguYll0Bq4enxnoqXSPK
D4uGG62HRPa/zUUPSJzDD3f1Lc251fjVXBTTWdI4+jWpR46haGvHPwiZtlUTdvISPQe83jRZSXoP
bo1KNZpSSdc3zlBfWbd62FKZKiDGCQEcUZRRR++L1PdPwxPu9nDEBrkXuGPsKTB6bfikdEqBTvjq
jOQQVrqZF6wS118WCMTPs0Qa+BPFDnPMyWDbe8tPsZGKgpVFEoat9skOuJVGerTm3nlZFnzM/dWE
lskrHvP5LvIWQsCGyq6XehhBkIO+dQtBH/zGfPWeFPO2cdv++nXjVNLBz256cV15smuZFGnSGZtS
KCx3jOpc4FKf5SNZi0QnMRTxn1PcxJZn286NDemt5Kx3dO27q51dw2X89u9475njgLsmowyclB5P
9vDC+bVe4gh37LKRFVw1cwfp+kK35Inmc79K+Q3uJfXb0rlCNhT52aBWoa+1TSRoLjnik38zrUnL
gsI8/GvLNaIbMGcbM6XBtLSbaDy5tJIJdwt3XRuGDwwY5odDUN66EFHgXrvd4cKy22SE9P/UwnCn
YVZD+o+w41tBUAYiMlWM3lEoTwrn5GOlL2bJIn8gERlfmF3/wCcisjaXmTITuQWpTIaPUAzBSkYs
BP5aNW6lxIhsRm6TS5Y8Jk3LKDID/EXSdhZQesLBuOagkjzyKEKb9tCUE7klNgaUTVTctG2pyv2u
2TZYa3oOoozZCJkrvI1EXTmOMC+Cgj6frJTwXYqHHjTPDSK5bRUKZnWCfrdXoVCGZ5k0cT2VSHrB
qIsbsE8haq5BFocmD98lnUtUFCgZ5Ht6L7VRxYJudxNq4rsY3rxlspH8cKnlZh/Kl9/YNee67sxa
kWXAN3kmARy+ASdslVJeE5kats8Z31pYHGOH2eD50g30EKjxEt3WcmrdokBy4TGiv1u7VVSZq6hv
DJ3T7sqF+zPYgQWThndAGKd1Y52Q/iZcw0b1EIG4yWNDrgy8CTw4ehg9mrZmw3tl/y04fzp1uU9Y
4kotWwaM7+wfF/v7rHKYSDNl3ENyX/WCdUQmVaIJkz7XHKepXvim4UsxmMI1RdR6x6BpRqHkvJif
7lZ7u5hYgQ+qaHpA9Cie1EMuU6K4uku1p+Mhr83vlItT4WXmil14O7q5T62Lo9keo4XRgxEh2sp9
y/yfcKzdjycsfgVuRAZQFbZ+iHDplIbFKNV6WSuLT7wT/uCgOAqfDXZBK1VAInCeAH66e36aPGnj
dxJLAIh47HQJcihVSJArPqtJeWWYx/AAypK68gow6om/JyLP3QDKWFn9pAr66HTiVskWmyn0Fdrc
gqRU0LMUWcc3krkJjv1HQFkZutSw6hItJAYtOeIVVo7NO6dheKvsX1NfZ4VtMVS61snq15dtOnnu
gr8o9BQ8Jmw1ySR2w54VePDg8s8tUBySTXWkIE1MuAHwP2zyumGvwgQhiAF06S0ywTeEOqOA+eg/
+jdBSZ1Ol4OjbGHoD3mIuJeLzdEmTvTY2JKxf1m9RpKI4lPUX2hIrSy4OHX+IJXiJn/d4D0+JJDe
HrGQQGddj9O5BIa31yPWbuMa9sUOI7QBi7lfJd0LD+nhzexLpH6DujlVfw3pfAa9dNbKda8dksaR
cUsQGTcRhd70TQ5M8Ip9ehapiR3IaZgGzWrRdjDgQHsytUxV5SxAYjWL6jlFt3LYevVkQsZqe9QW
ffujOhG321cCYadirHFtQ0w/9Gnwi6mMSPY/TPvg8c7kTM10WrNUBSPpoP6pFJJMTt1HNphZTxpf
f1Knw9Qo86WIvYfvBQONmUbzz6/vZGDrNA8+V6Ahfaelpf9ZwB550A5knlgRC4+NSht8MtatUWpq
zAf6SQ/0wHNX3ntSV2PwhNvwd65RO0wPuB2WI0kYSRqJXGQKctzb3QmFcbWKJBtP+QW58AL+SLVk
/5NaHt6px3Z9TEgscwRDOuWoE/+Z6GUY1Y+fYMfU9chbll5NNoHIfADYIkyaSPOqvoXUKmFw3Zsp
kz7W+q7dXe8orXvcy1WT6yA1WwxhHIseLpNtwF8HwmsLfHfCLE2+Q7Wam3xsaoMH8ju6McgAZDnS
Hv+SjjCWRItO2KH0+/HwxdBp6mGplW+Ovt7UhVC7hEEfygS1HKpUA7Egr+FXT4eet11H9m3fHAnX
ZE628Rxgtgip3c0AEcvhKAwgxSW1Bxgcym8j9kOyN1CRdaHX6X+zRodmLKtM1pudNqM9EKJ+1XyO
siCTdcEhyzTCvb6xNLs7wiXE2kC8Y/nBpAh9a9K8sl21i4KXsgmTAcV/nl7GkUztLVzmh7X9BuKS
34DFBULuQrG22Fd0eoVHk5MA0oTGIr/IdOa8NjLUwfWRWpQmEwDaZsoiIC+v7SI0gbxl5UWLN588
HNzesPiON8a8KqfZBM6D1Tpr/g2yRpKGaQHriQ5PoBgaHNyytEKh6wMQyzsAGfixoVJ6CSAKm5gl
D62lCKmsFWU/pMnB9dIebT0c50WHx+QVYfAXHaEDb3Sk+SgvN9GdXVWF0QLilzTevd5ZIQlD1CKz
O/7EGbU7uH+YVOW5WTJlNVZq7eApYdRMy+cnaWpyLxxXUVfy1mOLoZFvvPz7eAhraFqkmD+PgQjn
3u2lkXQsMsvXRgJmdXnf4gLei3cV+Q9Pu4xaVoRywcM7OqlV+/fHGVcCgrrcvxCFcHy99pF61h1Q
tAFwScFhC9CE5Lp+ZV/5UkMR4j7/Jc3rbV7LzPm2RaXsPRoiqoeVWP+M5nNFXiOqQnUPFm9r0k8X
tr0Q6gFF5DCGcw+IiFKcyvEH4GU50v5I+wHNNNazcEHunZilP+lHJ4SvXEckjC3Msyanc5IVV+pe
GDYz8xC1edC20hNrL0h/mjz4HNqCll5IoYQMXEqjjcbKcK7MZUDM5lHQItBHUCAcVWTAYUI71j16
yEyKSzX7wLT7m4RMw3frDOssIP2YxAbBmHygQBlAFJu8cgk4LSTbhdHL//e+u5Km8PH4JltV/c2s
7XT3n5ukXnZUkZ8PH2j2mRY0PeWvHuUXhL7mfg6LgeBRy6BT3RKkgw7eK31zYY+w45lIwoX4LQ8I
tdeMz/mRORnoi5y7a6xinfrT4yOE1eWUkGvNZ70zrm3+5KQtnnXGGBngwth2AskK4X6hNvhzL5NN
m4EcQTwXAIWKDZ2ckPby0YWrrprtW2G2bzbgX+Ycq7Ll9vaSDkQI+wiiDjaXtYEvlrtqCH5gMPqj
l40uolh+egC6GonoAp9+MR/idQpOB6CozYi9Txywk/q2WoO6shhhHrACe440N5wRUucnNSKO7i7J
CF5Zp5rpTWRjnyIy7yGTNDxxS/d7UnAJLswnnNVKt6kB8q2V6rUzdsFSFKmFj2gGXLhOiZwbXOsu
pAmwFrYaiyDbyiueL+q7o99OtbaymP6/nZQH2KCfPEtZnNUMRWS0YQuKQzk7WVCyNAvM8ftKAPKt
95BgdktzleMP5o4QE8rjuCYT9XSo11JlvyL/71GzbVbNf9D574LuX10aU8++2RVB8J5d+lbdYhx2
abrnS/9RksjPOzFJgUWjuka2bQrADtE2y7kWqYKfuhNqYpcF2XGIzvOjJ4wjv/0BvFyI0pRkerav
LIg4Gz41ChSX7Yzf7PnXpANfKlCLF0hwZrzsq6WrAypNDvWIpMTnDjVvdJf4fmYQ3RKiSE+bQuQ8
M1hDJjfYxJHV+WuopWUahw0ryp03wqpna0vxP1QbOJoIrx+goIfCY0jcqNZEnmyCjwmcI1RN3cbB
960FG6ec58d5u3t9Cj5aJPZa1kNY03/00mywk6/+JyF//ivwQa5iIckzPwskb4uoGGrtt4rDCbQ0
IOn4RAaFDhocMfq/wpX5ClbCkL0igYCY/rHEaSyDVXUgGe2LVMvdXaXKvhpfrRX2/eTjoXVIlkAU
Xrklnho7VpMvu3L5U38DdcP+xuTaxKx6F7weJryQLoGgYgoyanEYp5V0TFP9ZnibrjOKc02rOet7
5KJXZuGQ1Rrn85Ap0ZOUWiMFLuIiNVC+/LgOWUaYGMiWWAOITIurzn2TdwmGpa1Qa1QNfmbjbBzH
+nTjBb1YsLBjwZmdWE61lOYZI8MI+DAn68LOk5O7ljBHfR8mwQCz7KIKwtmV/KdhMakq/vLT6mZH
b+ozqW1I42CjmP+V72ND0GWeWxyv8ZrLB5sQtPvtanDjEsL6bBmIi2TzfZB3/3vA9Hr0T2I/e8nk
59pbDZrOxNnz/XhMNdBkfvTaNa7+mElmygqBSpWMJcReJIN3bR+pAq8LHY+NwK73t5g+e3+3CUBU
2eR78NDRC0XUPEZ6PY++pVwYfrBapJ0XpKKxdcOhDfElQxWJ2bNridt+E1JDM4KsaNIpV7t7sirp
hJTeOAjOPZHRTHWEm4dYEvLrmbfDRCa4S/fqoL2vQ5aic80Ni3Teighr4NmEn3C/UGjuELkX1IaN
ZeaASrGdqHizJ4a71OKsVhvWylTS/j2bFX+sWc6OlYnCCL5GX/c3xxQJXXsXbSbroWpeEgDJMMpp
yIQW3AJNbH7g2U1dj88dhQP5SDYzboNAcJ8ZfbhFmZfLVWpUCKXHpOkW/FqTbH3hLYfViSKzA/s9
DduAiS1OJP2T/chkCSsPdwNi4nfBdICQeLVP9x/XZ9azN0Ymf3nhBTnbp3rjYoRZYMnjbzDJryp2
lJp2+/opOmV6fU6TcHrAwrOOi6tqwkvSlVSgf3vyngiHcS5j6Iub6PznSQ0ddY+DBe3JvWYBe/r6
TSW+bNVWjzdzaxKw266A7wxiag23L3gS34DGBPVfojQQfRa7j2wS4Owk9vjGDfMwgFycNn0vhDzu
ecx/n+JBYc2KIM0345t59K0zEQFflci/ImSla4vDXqm7cIyeZhssjQQXMUBKTQlA/enx/KeEGn1m
405tNBxY8OcdFbt/wOTakBBfPbG6O+KMrdK8us4sh1H9euAYEZdlD+b7psXtivyyF+SOGifICMEh
zDyCrNAVssmqPLrgRSdFLk94Ko66BYw+zEhwU3R4OnTarC53Va9UHepu8NifDfno7U3Uo2liRYig
iykAxrNJX60+xO1eEgjc9BZMODgKTawtyNyZLWEwOS0yHMA/WSTaK5+HW8mgfwdO5MBFmc8QQa05
u13mdYXwTDNBZzYLgb0FBd4m+4+nbNr1vbSZZ3bHegDa6h4VjjunUlE+UfRjqgJv0CkmyyUGqR8g
adT7A56DP55Nn60eNOAQlWDevJNtOt2QC34H6gHA0W/ThoZJw8lU+hk4pl3hWkUFMHnhAhcOSU2T
3abg3C/7xjrxHU4oi0xWX9P/pk8SH7yG3jqaK3AVa7pjm9TEHcz82mKzV9oBVOZL2sXmK0lyB5Fv
9sLKWlSqUdYDbQ+pQb7fPJLtRZNkF8V4etajagHbfTn6eGC8zd0zu2irTTN6HISiwTGRxNlzekiS
XA5OLzp2JwQRnGHTLezWHh6waDQZcNMahQEXAoWNc0OXochKCjwO3e6mhmxYopSUhoDhx2rP8K3G
VUJ4SKKOTZblhXIZ+6K5tHWpWvPhNPpGJbNICqnTFjXtVc2DGRvEz6zGf6r+w0d0xIzgzvgdmqyv
luQmChDb8PguLrrpLSib1h7W1VZ12MMXZDF4YPN9d9PapXODP0koIuvvWw8zq5/UhnNAK5zr4IxN
O07/TZ0BSkxL4yaXcoxfsS+Eu6y0Ql8nk04vpJGsFBBt/9GaJIKZ8KKChT9QIoNiy1T3Xkn1rKH9
ZU7kFc+VwPL8vHz2vovPliEDPxjBT4yEIFJ6uHCV4E+c7GqPuqhgotCwQ4bxvPtX7WBXW/cMn+d3
kZrZPXp+lLiJNksSzbvCt7xCGnkdDBid/YbtTobH5NGfIuNNdM4CTQOzoMNceQdn0yLvyW+GbRhh
t7FpBTfLtHje/+iY93z1akK00OaziHB5D/O5wUZSZmsiJH4j3JMQFTrsmqkdKHKiWTnJzk1fr0Rn
FBoYGVY3KVZSWdCUe/WFP1t/EyFVCVXezTio+PlvyONi5tVDJeb4LqBQOXpWJ1jdnGxYmLKB7fG8
2o5hDK2kofFJxQ9nZyrBT7YBneU3OL89MGrX+1uQBE36qKYzdywjyXwgimtpr8zrw/spQhq/d07z
rV9Hnqaoyfl0G7RjWVZMKL0/SE2Udi5jeel6rIVw5UuIN5BJYKSN0aRoXRUB94YqpW1PK9Prj1x0
S7Ego2ZPPYKjajmR1zNA1NX68uy4K+el0npSBOPPjDAo1A/FuXVj1EUg6XYZWWrkZKG2Qq/8Z1VY
99j08m5qYZ4l05hp5XDoOYUpExh3gOM9u8Nw8ejQZBgwl06QchdiZtTmWzAxY0KsFssieveHAfZw
CN3/NhowqPp6IFyrHQnoSMW4EtY5XkqONusmys/Nxt4/16aR/pdT4vqUI2Mvq+QWAwUEVzDS9jEQ
Vl/Mt7s8ziVf073j2+PcMs0pWoOOk+Hh9ql5ZR4BNGqND1UNKyEyLdpUDVCMG63Vt4in8X1IlVtE
IOcPXOeFsJrq7uYCaErBLfWua8dHGg+ubdr64FeFw4me/3flFT/l0KeL7ET2K0WbodJy2q+TnPfs
X98BYqf/vJbsrspElI64ii74x8kvLyW6n8qsvBQcwRsLG54REAAC0IsT8ZaNiy2zyM0izJxhAexg
2Xoe2V0+Ni0PIciSauf4Q3WSgCdGeJKz8qiONIzrtnn7KMvyiKa/NNFfl6xXl5NPHviV712I6LGN
6NbkRNnw0W1P3fb73U82dHALHNFpo6oiPTyK/nykgeJQN3ZRIyN3uk3cl4ngqAetcJliAD41LwRo
nz5cfUWdBkbCdDPssp4Rs7QwP5IEswah4DwPjlIDmaVqptTTD6nSrCkgTR4+ZS95FkVZQ6nbcHjL
yVbLb46g15w5/JgWoSQSI4ofgbs1g/UFYL7XvucCLRlhNE/tz9EB5oZOw3pbFLvZmdyhR2/Rlxdx
Hoz9ne76+tQ8HGw1tjrA5kZT3gtgUZ4BxyqRRLfAzFXiFY2Ft8k2GRujDDDVWbOe/mUNRiwwdADY
2nAoiZOpeSjDjT/wpEOkmGIioIjz5WD+m8A1w2g1zG2VWPRlc9vjm7NtEGDEt5/V4vrN56VI13nI
O/gy16cO6/Rs05l+6TBNB8XKLmBXESYu6fqQvmsc8FxBkwwJSZyNqo3/8477bApFNro9w0xFyCB6
N3BNkJOeWY79WcIgohup94rTQb/d1ibzMbURq24XQxjm+JV6KkpKN2gTgdVn2H4HGvMIxEkCt0RD
U58mg9HMDLKyOHvvrBirsemnOmCaEjIGXYi4L4xe6afodCw/1ZXzigNtoToKpFNgm9VurGEuk/pl
7kihrZMke8DbwxgFz+FpQWqN1IryW8LmUf14b0zcaCfDgOKt0XaCSbFeQPFOJ7SxIOVT2JQMLiMk
YRGWfmcj2Tx2NQNslLIcl5okDhZ3jFncBshlJ674DTJMvsXJ+YW0qHxjIxma8mMlipLqwW60M4+P
Clrdwj6Qt+jcQGVcT/naJ5YDQn8G8tJr3kGuIp6eK7ZAFBg+uFu6T/b9WD4m9sYap71VzqCKiUTw
isuCdzJ+FWqtk2dO+r4LCnTFvtdjdtGxldoW+SLc/AQmhQUDiWTCfsc4POg174IBB4On9N2U8BfR
FBrb5unsgy8ZhQGuH+FTw4ZwgDbonIRFSXLV7NvZy/zUl1imEsbYdhWGOAzQZ5bgNVX+1kra3u9E
YuYFJeIJOyn2CRTa8Gr83jzbgU5IzxFDLXitqq00bKhBjQMbO9z/GTIAHGuiyT4NEts2BYdm9xzF
UzwQsQHehb6i/C3xpTGGn1/q7BG9mXQGbQ+CGqdok4TDfG2yNV3iBjLL2vz5qHgSU+QbSQRQ0xLk
YsvrabipnEC4VLyTnWVSE04IiESExhovl65j5q7zmJsXySYc9pea3EaY14WAGEexxr3jqSxaAnbN
NcsVSKifFNi+nVouHpOtis8ylcVbuMqiq8DVaQ54SxpZIyrgta7s//yxgUzhKFqgCwtI0dapDreM
m2HsAbB9i2ynxLBgxxORX6infBTcj6aQ2GFFP0Msle+UcGM+TrSA6I3ScLoGGUF0AC0Badw2poHj
27y6Un3zDOu0lne/g+GLVB4u2WlQ5P/rHCSlfwMzXquMWPvcaH5PAbBCSS48s2I8Sc5iIoa4wivG
cjJ8FrW7AfeI7oPONr/wDL1IaPGNvVeMRZp0LRNahE+eZ2mRAZ5teK5A+8ze232vHuv9wuFz7KPB
TqKhsD1u7froJg7N9LyjUfijsjGqmoFpxWj65vt2npXuCAW1Gr+OhoCPBIni3bZpdZefIKU0Pdyk
zPfGuyVESrxLc5hLxhx7qKmQ4K0g3IPA1nmB8JV7gIwQOJ2hBfk0KCOu71YAHXO5rCWWRARqa687
rL68Or7wmD2aO0zb0IdEruyAcrFT8d/QdLGvR+TgXqsC9fpzGcsstXaO7p1r8lG2PNUoxjRqS8bk
5xSdpKPFvm0+c2qrhsXYbriN/Y/94mXhwhUZeSFyo0BEn7ZzFgcgRf8b8FXEXoSqNoGkE/3VUbj1
7QQMrM79HOOQcmJtykn27blChQ6hS3zQLSHvuQGTgJPD+suklm5QYQNJS82a0hTwVhvA2cvIRKFE
Zypyktzg86YdisFY+Q8D9KdjHYswNGXs4/3jw+Nl4JjiPK/2UowPeJTGwhS0odrjb+jRTW1kUwbr
8qx8ucyDF18D3/XVX7sDmAW4QyWu+QE7JRyo7KkYOFwk5pzR5oGi4rhE1nqcp9ptostT5IjCMyIs
178whmKaVa5xs7QlyvAyf7xqZXRCamUvczOAoi7b/J318Cs9U9r5MO84sbChssiVs/fA8AQ0s/rf
Gr7VXM6LlAZ+UOeDc2doAqjORU0Le3Ned/Y2VCa/wlySBZ0QFV21rPoYbcYd8GdfGWDPS18Y96ve
DMRrSBXgLV2Ztf5pk59/dMgY4fikMwTF8nPUsqjs5ZXIdULx4ilbZql/rRAWESRGqf4gCId4LOWV
GSP4BR2BRNVVmRIcHRB8jaCYQBgHf+4vjA/xeKFTb7IrmrF+x9ikYlI75b7SAburamLT8YJFHCDD
Jhh9UDbC9UqK5ks8ILwOJfavUORoI0TuPsbjBP6WFYiWQrL+3rD8FViL/L0tYsJMnIIa0CEz79/b
mNgwueIOrkUCVvRbG36qNTz2QzjP9WnyXXqCXBgaiPBvUoMRP71HqNkiwssdDfO9PrPMoVN3Q70y
khhXijuS9i+iRdChFN7sHAqBybCHRnzWYCXEDKAXtQyd5rnGQR7RuzCXy5ksYnVa3S0yf/nphBKu
IKTbmAkRZyX++jKyhxM436tMBcixuy/oovXf3vg6roIUVm3vT8SawpxEnO3FeN0FLGrciTiQLvnz
5VEBCQ5Ivyf7XIMO8ctZne8n3MbJp+BEe1zWJ4fYSvYxA1+GQx26xMndKZ/XT8g+apnwc0w3LoPC
qxfDTkDJuHooRcPeSBD8XWC4A3POorDnpPhaAxR4wu3k51FpJGtJD7DTpfhl1P4t5XsNAAEjwYNV
b3qx5IWNuYcYFE2ODgqrB1ipUhodcpyhXeznZkoOt5QTqz1G/hTbkKrSv94w2CqRveZIQmO+Ao+V
hbwZ4d46OWHdC/odZalPCm3VhY+cREYXb/17nc9xvkFc1z9AdAJBEOOpIZG2Gl/mFR4UcFs7ZiVr
r1tTtqh1swquU1UqdggzZYxXFkLVm1gFm+2KoZF/gi4npAuVvtZvzOi3DPBsR6Vj3+gC2YPPepkE
jxtLZJ1jh4HwnIV55fxqrJPZ33fcHzlSU4JvzwMvEox6ybHYuVYYIPznBAO4bwhLQ/I+XqPGiQ10
4+K5DEMtRSQrhFkI1OgOQ+GUV5iABYQ9rOSoIu8PdUcZvEjvLc7sfZi/AwtEJkhg5hpLhVGgsx+r
yCJesHga8SFhWp4XBkWWdEYkKMvxr3O2ZjrrPE/zvOQTPi6fOw1Sm/S9/vNiN4wG0PmEZp4THiJi
vkGDstcivhaFO+yZ1mCk0ak+4g2i6jK8TiVrLyG0odIBiRz9AJ8RQlM+QQk7r6MPkBlo3aRQqbFk
5wQcfl0oWa5W657XoFjBZO2sI87TEpv1x/FCS6vLpcSwBvl2eAh6PLEjbasGyGaYMFXXvduWd2Qa
ZES3XAoW3UTVhCBARap6hdkc75NK491UmRFjKA7F5kfODX28+v0u4L181r26BxukZ9+/lOOzDriX
XFYRETqVQVE0RdWzUNUlJsGFzMp/RkZ/ZKimaBL35+DbpfzQv3daEBTRj7H02O5VAEVE9S8SqmtW
RLnKBil3C9VEYaqPPGnwiuH0luWoMgrshKk0/GnqpJn6fse7f6wIFYX4CD+01lKtj1VzGMZbheM9
6mo7QKfvkWJ5UxL3+qoDczaC0XVL55GenFkR3N1IlYUQwoDsiyZB8ANL96MKkgCTVO3QI8bLUar7
c3HTUFa5X/s1VjTK68hcChDvha5Z0gea08owWkdkJuVG+iN9DaqKy79T+JktjJZ1uzhB7ufQZYUr
CY0u0eWMrVY1SPc1cJvnpWXaK6ECiAZ4MrDnc9o5FfTj9zTmrAq/2B2MXLbSlICR3sKBqrFVRmmP
/5lljavZsojjE+tnVPf1EnMbYMCAYt75PryHhmymK1nyiQG81xcCGrednln8kg71svnbuhdw4PQp
Ch0/mZvKNgjEtNc1b/CwjNn66qv4lTO/VzUYAZjzXLeviRxNl1/52r4+1k3zfhhombakNxgTcT5Y
x5++jOZL40xHiCNRQ9woa2aaNNOOM/vkI7menrXCxgWr2oo816HiES1CT+PMwuR4gI+/j5mpp5iy
k9oZkIJIQ6RIOQ74mAuc+pOZsk8917ApLiDhz5ocsbNPSVdgCak8S5dV7vtaF2iO2sXGaanEwWve
BKyGglnS3TNEe46153eiW6V5o+597QjEq7coBeRRlD089HjaoCvGPdAGPHnFG29hJrjBYJYZuWBG
0/YMbiJDcvWa+EdEhhmSGFIMwYOUVN4JoutbUBInc175jTndymxPFjlqHSk0LnhRCyGf126F5cuc
pyuEa6eC9ukkKKbG3TJuWYrMN9Ze4xIGB4fGwotEXN8GS8tF4jUjWX1B0bivz1PCBLvOJEJz/ghx
m3/ibGbCOHmXM/7tTKEsGLsV2jai0HsvT9tqhM/+VRDGqWYRMdJ02GNGAMPJvg9pbNXkFkM/o/Yq
ibKrgL5xJzgTRREWnQXYZTZbaV13oLXA9QeiP0gPRbjGOC/U8WD/WBew/dPLX2a5lSdkWOaVJTdB
A0MczuSXCOXm1vvW6h7GlfSAqoJu+zpwA+t6OUD7THrkC21oQiXyUxzUjtj8QC8BURi7Glwnk9Jt
VcTQb3aGMgOVpkv5KptQPqAu5NbT3xLLO0/7hwkbfkKtxdSwxYlnLJ320fWxuIYsGp2Lpy58yVEr
4dvF9Fb/CQcgGQwRvObawv9B0r19kO11bdZJKv3HvMuz3cRYJ7p+/6elKvU9H+8y37p/Cik6R7hi
n+7N8876UHp7KDcb2V8aPHw+qSbb73Q+eQcu+HX/739hnsb5DHsXhmMNkeijPkggLJm0Mo4Kw/Ui
BvOZWmIzJsAAVOPM1DPCsEdPrkhmKvSY/tMrdx7aPSv9Q4wmmuhUFD8vjKCr/goDZ3GOG7R/myJA
WdS6nIrKHwFuGv3/HPoj7tb1y+l3F9TAS5gAbjosAOzIgM8THmXv4NtsHUWbaJMLLNlshJv5tYDh
zfuLREdhmuQO1rla7LTF/3Ds8Iz3pOi+sLCWMLllbWVzRkN/yfcPCAvYW9Tk9cStHpfJT2WC44Ai
kMQz9lZU/Tw/20hH0er8vvXqkaMxuYJO9uU2Gzho7IyDJMsdBtCsQa4SU4kQR88NP0T6SeEPArad
yqbWKd1MXrRACYzEJXHbAcm6Kx2gSdI60fGbfsPC7sgoSmvEcD2HuXIKanriMkJS05HQhq3RwPOW
DA05ZrDl1sx4NhmGvEGht7kFfOxAXxWrhnViWERLpzSCTB8rq0z0eOzwtz9s6oSKDaB4YyUh3FZJ
B0NoAuKmSPB09qXPsWGtjz0BIn4VFI6jujnDcdNUjzjchkuM1Aq43Ca26OTGT0h05p8cZbTEVuNR
jqunMKKr34NmGHOMHOZDZ+v1DIf9yiNKOui55OMJDSuJGUCBCATUwqYxDHeZLkVgJ9TIdssNeBn2
gHhFObnFf4aVo2ny8A4z78g07WDyPpikvlgxARBrJcxlmfFKrTDUO9GJdQu63ndWCEXdHTL3OHfT
DuUyoO4kcMx+USljdtOXeLAze1lR46mB1DML7eia6qKuUxl9qGW8eumkIdX5X9wn+JHw9jESW2uX
dNodqidDfDZFvd0qqpBn7RIyQEcn7TF6zxef48LuyQcVIbqfeYwYNgGZvAYcGJExo9/Z3ZLWJBOd
RsSHKG2r0wsxwSwuugsvpJiwjRYxIe7dLKpO9XO76A+wuAq/aECKB4SymINVf7A9mJ6c55/LKhdZ
4rWPlPghNb2bSYE98IJry+ZR+i8xECHVozA1lr3V+Rw48adsf6MJZQram3emRWH9jlt0o9SMzPRN
uBEduL+lk2gRi8JfrvjVkx3jPxMxrEbPAHAZsxqfPXS+44m8BYOliugy15HQtGnt5F71fubqhPM1
BA48vlK5tz5+0i+orr+q58qKCGjAIvqbxbg0yOLIYlJ3ypNSBht4dbAznrF8e+aLz0UoL5B/c0m+
HUh9L2wXu2U1TVJQETPLdXyjogpaHgEdMDAzrp4SGoOLlVFVswGGw9aOdPf59xsu2fkCkF8kXsYz
0Phw3oi/qRFQPgqEIcnS+Qf58dUkAo3FeLKLpYvOJDqpxnxmt6RcN50mHunU/2SsZVpAZTjGHl2y
pt4UM0ErEwrDKcCnWkzpIRD20HZbrTuDzwJgCcZQJxMOaRWW56fl1bk/KrVXEgb09FnaYxhYehS3
RDVaqusqb4xsRlnkE1p+IokAj8IO8HLbxigMU6hWgw/bUM4G9g33oyWD2JiaxtCiTbRRQfdQW9DS
WGEo1xZi7eaSlkO/MLfFtPptT3kmS3nn7WAmhPcnzjVpgRyu/K5r47VB+cDAY9sj+6t54XTSPRLR
vTQIo7iaulN56NBkaHKe0u67oaJj8WjqPeWYp7IBUjzDYMo2/ypjV5tq/j3kxiGNdk4oIbQ9f3Vx
/gPNPO3bEK9VMOeguSv0F/YWd5jcpcTk6bD1xehTwE2ZFOv7Y+QAFbUmdGHIAllaV/b0VLIZMYWs
gz/2UkTF8j5zB4J6/qd2JEYYDmsg2/DFI8Vo6PCz9cayeKE0bTEEhf0g2MlxxiDuoLd78Es/hUiA
sKT59WSuJ3+4C3fAXpfCsQCU8w2YX1i9wq2ohht2OQ1FV67fjRc4GVgLAS5xyZgXS4eN6w/8IJ/Y
pMa/yUzjSb06EQGtI8ozKeFy2oCBHikDVyrN//Du/SS30bm5XJFJU6MBAgLhoAJ4j/WuFyBzcULI
GF/5/2hlHxRQIJvymCcA4ZeHhb9BeXCqqDP4FwVZFs9AyXfez9akDAjevFqDHxJ+o9wu0bnPPCPB
lEXRIqF+N8C4im6DqAT6iBmzPK/L0r6FRSpD4IR3fZrNufFouazvhJq3SxRRyKu3oT6Vkrmdjc08
HXuSXrgKpY3Fpfu/Z0w/2cti5yQfZ4zI1hXTI5Bbsfv+TThj/JPF77vQommFbt3vquhnPzs1PQcQ
FWStUQZuMvuDX0DemsOCmTe9WXP4vL6qVBjt9icMfHE/Z9om8AJwUZyAHswrFVB5dOOTqBaxmhOG
Pm3eqKWO5ZfTIj+T9/zs5s5NMQ1d8ryck2LJoqVEeq53TNkqUadW63gXmSy2Lzt39EmBuY2tPnlQ
rNXpLZm/zMcHDwgUrwPT2O6w5Zg1Ojf12WmXUdCtwFQb7z9IUfte8gvnwxfUxTUPEG4OqUzHZ7GP
kmsq2xdPcHj2ThrguhKYm88pXDLnbgHwmz+nI87Tz/+LmJdOFk52goRImC0WK0BiyJUyzeIJmjFJ
/f2y7f1Kd+oTZjxgD1qLcrbFNOb9PhTi3avB0xuTJ7Rpc657pOnRaxZruHvms8S6b9P7gZLoRk++
jx1I6wan5x+lfu9U7HpmIt7fr/0wuAeqBYKTB5xUopreI1EFdm8MyLv0BdzWatBZyGtlktu6Si+d
9pMKVGIu6KyPSVgwbvOCqF85i9euXeI/TAXC9pMWZqW5j/RskuF5BECaXSZoODDOocGj2hZDmBvk
ZGJVST1fhcxTQ40cTxfjDzQZ69DbscrEWVtPrfDZrhVyiVl+yXUUyb3Cwkt0hfoDrx7tDWP/1NnU
8tXM7BCQv/HD8XGsIdPGVBHTud0bzUA2KSTUlTPOP8e5zrLBE50vgeFcMhby04PdWJSIfwzFwql4
t37Mj2ScqCrREyDulbixW1Tc458j22gffMirQLiPVZhBsWqmHAvXaxU5oQ+vejUhCsfBuiiDi+04
WiscOZPGnod7YnEwWfGiDGuybJtLzgan61MXBrSwav+JikEsE8apAgmm0XP6tTOs0ALgqOGIRTJC
ZKar/omEQnjiUEzFgsa2sylpBIVQCJ0I1Krg/ZQrAn1sWsSLM4fnBHiKosDNm9EjC0eq7vhGQfaO
AdmUb72NW0u5/EhfIz6zk80QbFqT9DAZ2b9+YNSMdDfXZmeJbgR9YkxYA/1uu2LUwuAvTe0aJOPE
8qf8CYdN4qslit7yYBTqx3oAKEIUhRz8pqPRaug62tNtRAZ5trwp6CR2ursis8MYD70NM6Om04kL
gaVG9n3xOUjTjntuf0gOxa57Cte0u0jEGvgl8TDAOmd52nl68u5TRk2+PuCElzzji888vHUEuZ5g
VJaqkXhkWChoBmFU71S6+oszJKCTFJL+lL2ZAFDG4ew/dDBMqOnQ6xDyieoGb9Wx8iffRts5aZnK
5I1y/1LlnlHnRTwfAISn3jaU7rd9iLfpI7mR6klz/1ksOsqfgTGblFDLATdFWrk7ny6jd1M/EpQg
Adb8OVWYz2ygl18Vk5guAzjIiVv3BaFYBOyBjyoZPU9TqMWM905Q7PRwIaB/L8hJQIZV9XBr5sND
rGzh5e2i+x4xyP5t17wTtPaLrNc+QvJIR6Ttb+HuarbprYWvSu8HNuK95x+UEC3wU/6p9vHOqgpz
uYdfMNlb9iuy5hJw0tJmg8NlmObiNkPYS6t8OxNHKqOAlwWHR/zbwM+/JXzvhLBaHeElQJ/Xr5h0
vDuuzzF7BKZ+Ok+8PwWfzwTwiF4qy80IrST2fVWIDjMIQyvlTU7cO7EX+JvYBf7mvKYrvbNjmUoT
Nr8zKAob97+QKCBPOfyr+TNebcVbktSO8KELQjcNIlPFFXbh0l/zHKnfalg84vr1NfBs+TXra0hy
02sWpkAwS3JIi7jb9MQvxxOF33DppGCTcrsOyQNxwTt0kyDW9RZeTXbCSwrNEijgV9YM4vswUC4z
/NAuc5yLh3Wv5xUTIG1JloxKFk0PEFtl9TPB6ou1TCgSAjn9EF+NJBrKjfkXm7XsRlI01EubAjIT
qFLbIil0PBvHI9MvptuLUi55SjGSYr8OxZQg+R4tWpUMCn+E+GNpjGC38msW21Wv3Ha8Lmeo0Drp
MRZssD/+vN8RPv0nmPJNkymV+SPCX+acrreoSP3toBYaHhBuAmCmtnEc3LqgtKOp3lOYsKS7dHaE
PbKv0gB1bz5WgtTWvAhurbp6bMN+LXAyh3JV8FA57P/1a6yZYU2A/9f2XXWVqRkzFNKG+IdcPtZT
kIYvVycNUG3oC5QA3IT7zOeS3wUGVcqMejZxf+ziO7RVtGG9vGNLruY0YMDU7QnN5xy8dkwQQ9CU
WlGz3c7SilDJu+H1+RndHWqoBeHKDOJsO7OSvycrzlOCDO+uqXQWEVq9Oe2fkqEBF4JpkKTXXLt0
LTM56fqOjM0r8v2Nu9tT6YFWQY9I7xwYIZSfy+pB1nHSDwfODbCIgQaiY5d4t/3mf6BQmJcwNmuK
T8dsQ7Cp6ZSWOYO/vKgErsI3/U1Kqyj3PZLNwOiyTmEuD7Y+JHIAwUJ0u3/kwJ80dgLvUY81Cv2/
lIt3rtTixedxWrEyevzNUf2yv+CNJDXffhWsm4lf8tCkKPIsX7I3gbdwdRrX5faYo2sZyntp1eQS
L8/RsytcIBuJHESlEgBJ8hKzJIpul2v8w0yh9I130LRxvRU76d/1WTlRBnw9gHKckt+j8EKcxkEL
7gTd+IkHU3XxQsLQM9e1wqvYbtknDXn+Lba5puP0CdNgAF4/S2KpDnk5nzVxnrl//X175qK0QOFz
pjeHgqdKh+zCpGjokccjBH9YHUp5qO/DJpBr6Ac1XY+9CMLEX4zn6NrvH9rr4hGp78IFxrloDRco
/SnhPLygMsS4c61Yqp8BbOwgV0y0pzrasEcoV/HtyQmObS/iNRCnO9Uq5Za/ajqUvRdMsM1GbPNS
cH+rJDptFg9eeKm+46WaVJQYN/I2YggLJPkvMAaqTpLBtALchMXJVrGNPiK/TZAMaNTkKI8qXvha
RHwim8oSNRbDJeVhD28WVNVOgB0HG05CritGwo03D6/NihP6jQFX9gh58vPDlVjQit1HhQS2/tbb
+Ue1dpmMg34UyNLXolFx7Irc7EUdYOqHCKAw++BmmDmhJ488t284DKGC0+4PVam/IITvHS6Qo7ml
La8l5K5+dh9e+ZkoF9pfEjEje4Kdttctj3cXF+dPgMnYiZx8K/ClUSk4pF5N1aavp3bVMSb9xd7B
ZLr84Z0c0PU6YQpBhuV5VEWWK4FCAs8Wo8k7a1sf6fekt+yezKaWaRYZx/i81/Imj2eKlImMJ3xG
L/xTHXfnJyfuD1wdOYP2Att9OIgzk4mAN7KqheQvxqvjViUo1LdNr83yLtTOoDi/oLjqSjVfUmGY
8N2i300D1SLQegUMnsloTrG7t71NoGOvQo5gB9KBEkVNegSlgFVZuNAKv22Z53chN6/mK8rzfVDA
KyE7lcgni/ulZz/PcYTqis3G+LZ7UFDoNyuPycwdImOcDD7SoRVJH4vZMvKdbu9ltayuMjRuU8c8
bOcbM/opn8IagXA0dWXJU+609RLYpFcH2ng05xDiaX2EGqnDQnNRy0k+oePfq2r89PpUvNLrJAbY
DACoFDRACSXb8e/9VPGbZVhiEEY+R2BpDwgECLzXwjGwwuI10ydC0UtgrvG57yUO2onOcz4iND7F
HN4PYkVmBbp9LDuHtTU+7/JzwR7qrYLSWMZATHPvarRUiTwILHxeZesE1s19SB0feJRxk+v2mpmT
Y+psUSVgqWG3RQNyEycP+3vf0TqBw+Q6/g4EED0MINeC/wvRHttW882GNbIt4WSV03rxwS0aAYlD
/N92vZcMC/6MJzute2oQyCJHHpLcd+1VE4K8D04CCeaYYYoXxxrF9Quf41bALs944/5MLy1CY/CS
fiEGfYUFXka9EJoVSug3FAj2hcvB+V41ULvNshegrg6XnCtfzZcfD43yPQqDDrFCRb/Zy1vMaBlE
Psjr8Bfy6+o4Ywh1M3G/g20t3iO6ioz3mAyuFkbC0GhTKeiPmPGbkb4YXNsM+mUGgbf5lj3HPB3a
1uvYXf85ukJ2takMF+QhznwUPsvYmgNBKOty0e7oZGdva6pJlap8GNqgffRcDzzyEO9Ue0NX05F9
zHoTJCpelRsbJgENjSFTkm+nXmSnPuHQyy0y5YYLH4A7d8Gywdf6KN4lNkC3PJ6FZNSZ+2/PIDuU
49H9rLjo5d2Tq0Etl0U2Y5m233mGjDIzlzwZeRXSIsm7Ohj+102k/pQYWO4k/HrmCqbkWAfM+jwF
gu2Y1I84TBSPpj5SwZPjpMeA1QXYlB4nXmlXEEknKuGKclnkMKAaXmZ9cbWqJcEwUQuZzhNLz7Xd
AsOic+ntDCiWHD1vi262oyUEIaTakKy0TtwzsE1IxWZ1ZnDXc0d2EZ6kYy5FHkDsluilrdy/iHhG
wzvSJYJ8gs5Y7iS48ukCq2g+50E3NEvYJvxzCk9bbfcw9VaU2k1MQKwlTAXBkX6crbwRU1IS4jvc
AA203y8n9DMgCIBzAEe1MQeLUOf0ckpZe9uh4MPxpb9+OZhGJXFnfKAbPLp/kEhLbM4RK3xqTNZU
38/QsLTkEY/faqNQDehscyxaa7bOt+7R6FGKiNgLbXy/wcHrgTHqdTYrxUOxsfOpmFeakudz57fr
lOdOc5bpZnVd0LUBQJFJ6VQ0vPv1cSOJ+MVncVCbIp9rKFWbcuzwYd2Fgs+oVFxZexeDMb0YR9wv
ZKgPfFwA7syZUryT5TXaatjWWqOWQVdW6ZXaKXTO5DULfXTBeuzynbjFyH2JGYy7vocK0B06AMzq
SKKd71+Z+bXYgLxN4/2Il04rW3Yax8OVXZCMVTBTOnq39DsoPMTyyIrOdT10OGp6FNH2gGs8zyJz
uoRLzbYNrnf52rqO1c230IEtTzcpLIi0xa3Nm5QiFqYvJkL3sy1tBVNfErh5XyC/4zgrltE1egkG
1M0iqLT9nQ3FxUG9uQPSm/9DZ14Sgi7SHwLLt1P1WZoHXx6ugkwrNlS+b3LESBV7QMOMqQqMdzlr
EufFFR299ajc59cSDkEC5F/TJ20pGh43lcjcfNqozwExWmVxGJNwxc07+BSREBoX8tinJtkAmCUU
7n01EG4TdZ2mCM8GaosQeOCftBg46ikOc5k4t5rzYGvVWv93slqb6ad7DYaNzbxEg/+JuJXasfvq
7N38Ca2JIssnTxZ6jHkDt2Xi7A3Xw9BCE5vYJ90X/JLMrn0jmjFoPu3mVG4YPc8TBEwVxtaV0AsP
SpVgfygCB5ZEKIuEGwqyqKhg2JztZ5U6uW/Po8ZnuXgnIvZdFEqlvhiI+6uhNuaBC1VPoJ8EwA2p
RzpJUoLDQj9sAGLfGtVAHdw0S+LgkG75vBcjVYbSn1cHKHexR1F1XK9WDmeuNs+1XfBaXKGAOstg
EoFsZ4cz8jZYwYLdtBhYslngfXcETiw6GfLyaMiyToYr3bLzw0fG+oqPJ2De48LWBwsUMQd4p5iH
aM/AxaqsBHykJLA0ujtxW0AYDBPxbA0tckZg+Wfw/JWhkOM27wWhI0xrn/2oXmzbNKgKynkfp9jd
7/k7kIYIW0nFFy15qu2pSXXTqpao0QrT5nvercXruMKdasky/rha0mEBoX39Lt+FXC3sT9wBQeQ5
kc4W1HWens85wDcF0E9g6W9P5zy/SodP5dwuy1/H3felZ+NkJ5v+5BtnXSDPme4/4anhIzasiO5V
OeUk77GM59XFR/EIywb/6/1569MyvkpvjA6OG8O6NlhXQW9bdsaPi5PiLKXpXdkk9Lw1+r3RjM1Y
gCR6HBQQQel4q/nYaCJvR8SIgSHXtmii2oI3m11dK/knpGJMxCv2oKNmyAYVMVQ90IE+zF7n6ltR
sniz53TjGg6WqTSuMxgoL2AApJVL+h+CNs3223RC2Et32S23vY5rTnD4HbHm7JRQkDzQtPo9qkyP
EJ/CvIpJZCMa6kWjOHU3P3ZV0XsP0EEPt9Rsgc2UFFswT4PJmj2Axra8+qFoWUQWoZxzJIh41HFH
kJgKtYxJeOPB4bHLHMlQu72pX/PH44o7d+PuFnsRxOdoIXt6CJBpQ4yano7qTeogBK+taEaK76XI
KMJrOGUv2Db8FDsig2ZnHhiZD8yqUop6v7JyAaR+ZxY3mNdXpUQ15rdhI6fz/DEqe75LFhl1TB62
fOZC7J4PoEnvCVd9M5oBbXuB2WSPHwXsUNFdNAjZih3THIRUDrweqdwUku13JDsLp2FY91DdsaF2
VFbgjUDHT78jsWX6hYxtvkmkU/tFQ/ANjiEOn4Nm58ZII/j+tXboB5YyJrBlCwNVJRY3RuY5/W8H
oL9mXj1ezLHedJZsJWUB2nc2QvdUslZ8wqOGsOo16YbY28sYhqosxBM5Tz3/3JrY2LTIDkd8BL7E
DLR9PGQf9A7fVO0GF7/BH78z6cOKtEOlnSBDwG6oGnNWPKT8TEB00xpmKEwD75lbsfWNHndPa+jf
h5wILQyMzkoIdLpm0uVBw/k3MKH83w72lo5diyL2fShe3VB1PrcKuZ4WKYX3xHBY5e/Of2n7KplG
Xh4tagfVdJZ6nWMWOa1EZfV8MZtkZQpY+WOaGI6yzmovtUXVmzwf0TgJDwzmxASRKednbjTYH7jp
3KbsQGC2RdAxGiw8yGLqjVcy3J+XjCuHmW/F6z5yiqhz2GaY5DFYOxPnIUDEuiMfEwFRISqzoYsK
v6JZV0K8dqB4DZOdwO/NE4IKCJmVJWZUf7hNvZOnjfaLXEDYK965hJoT4DyEH32TSYK+apgj3hCq
GWM2aaeLimtKXulGhECkbTDLo99JhlIpV7FwKNMCcufgvwUzkBvDkiSvzjysuHLSHMr+CddmVEFg
g/widP78qujZQ95fFK5IXuN6K5RNqJEPj3ASUgw/JUnIRO5G0Qr5uuZDnwXblvWhpYXgiOQw28Ij
0aPnk2aBIttxgL1o766DY65QFeR5xyye+ktkILM6PHsX2jZ/UlPtUevLN1FHL/1IOFWm1VIUNBZg
rPh3LNEnq35JD3eKannCUkAqa59MkztgMz5pcSoxC1QeaZ0iIQT+/hh/lwnoEXKU/WMjhTBEpTZK
iBWyH6YPlmC/OLELK9lqlQve8RV0lcbOHKu1tDsYww4Eiy3gJGdvskS8yUbeqckcWgKxp7rvff+x
YjqvGWa1KSGXLCaV76zpTGXvvr7Ji7xV9Hsq4P3m+ad4g6yaVzxjZePb/DrgBb1cSW9b3H6zsc9g
YXllB+vA3S8dtHPEH9vqGL5L4E09RATkLzxVLBKFnt6IFGk+5s5KLYp78Gpg8b7m8TQCjRKA4JWb
SFV9KaqjWPn9nR/7p6FzDX5PPUYLx5q/hw9CMgHxJTLDvzYMpuaqX8CeaerGmFcOWrRHxp10DOzK
0U3pandvkrDFP+LD4V0ZB7wTQMyM3HgOJLyV5dHUxUGtSyo2XByD8Ls7IiG+bEL1C1CbhsocbX4A
Gyl4fSzYcu6E8+Tg/oQeaVwqIWCo/CbxvsqJEAbfqhik/vC62E00OdLS8M9w3mPw0nEWySYuPAio
A+y9gVqfyd9EuQzuwSRBf6uuTatTMYETvMs65GyrK8fmEzS+/6eiZfuiM4AVxp5s8KhEbYzeU/4n
1g09QEab2e8uvSfztpjcXTovOkURngvzuBWpSSk9F3XlomFfp4XqHneWgUdB9FQnC1G8wI9Jpb8/
czO1S24rbPUBgZHgftmYBxSlxuGlYj2pycTvrcrl0wX2VfXNA9ImJJeAkhoRNNorn9xYlz3/oWk5
+SJMTwA3GhAqV8mVfEtbysdI7ft+433gESlt9etl1VplMS4CfYfhZmHfEO1N5qOgdiHrl7M7o2TI
zOStrb18ZIrdnVZhDe9AjfV3MQG/wfnY2ZPvSb3BKgkWymfCvq/91tBsZO1mZSE1AIEmHDhHI8vo
ybADJQ2xZUA3/dB+X9dxwUhpgEOiCNL5Bz8qWSg3/gByjQyCgdoE9Dqk8vIJbs1Y+sutdTuqvsv+
4bu95zDNGziz8Kq4bIIF45+RMVgWI5eJLd++6vEZgMUDY1QLCBzb9IFCUU0UKCgcYDkoWTuImwfN
Tb1WhzpQWQI94wT6FIbAGo6pjE707XF8yLbxy3dIGQSVxHPQjxwfGbDsbxWorEGn6kGDCHpL4E89
QOUCro5Jbvl+zxaBWpJVQNNLMdIuCk4IjhVNIfpohcmwMGCMOMvUgi710EcrobTnvNaKk6VLt32L
amSTAf5hoQZsbO3HXglcb3gbOqi9A795xoQz7NkvPQdxL4Eig5NhTCpMU1WbNM88dasFYesIoNQP
D/GwbAhLHondXCdjmLS1xeRw1VzO3dggRd7xWnTWOSkB9Gwt4KfD5fNMAoPPW60bHZxR3iETY42c
curg8tq9EWKgKHLeKfMuw+8CZjGrOCo8Pu0s5t36WbXkL8OnFbvcuB1E12C5Eeauigpbltezuv+L
C9wOgt92VtKsT8UXWOKI8QfkNc89LPyc+chAUXPc07wWJHgwhj4SaUttw9H9M1rmWaGnXTP14tlz
Vh9JZtGjWF5TEQyndHro+5ZjOZs0ui+mGnLBOMMdSDK5fN1IHxLrugRb2IxC4nxs+jtGCJMNvtXT
Y+BBE44am62DwoB/QR8P04Osf5j1U51u+VWyrI1atWVrlHHBiQEofcr2iL/yo5d7g97Y/nNJP8Hp
InPyBC2AimfPc+ZE18A1gX3uDFfWHOKjCuQ+Pyp+Uw/P8Abjf1i0tFuz/+DrwXG1E98nCrKrY+P6
htz+sOM1Y7zS+y/2Bo/OVgzsFJlAoJ+p/CgF9JcEzD/StdgJ5LKc9Ebbjk9+Z7Aq4S1tsp/YdHdB
l+CoQSVyUNotufLWsoWLL+XNXbvufyejkR3olSu/M5dewO5cd9LqHrbHQllUzH0SDCkUhaX5wUeo
N8KkLYi/pA/p0zHktADAlpA3B4ubArdaYFrjtxFGFGNxWjMiWIcpTffVRZ8mDnsnasTzjMog+ti+
UUwbbDMnk/CWL+0AQpmii0WXIakvaWx8oAxFTBuYmWzOqEAhZ7VuOlneqwRCIcw42RnxMQWc7EQF
nZFAqftIsNopciiBIRTGP2Kvm1Lxc4lMlHkwWZkuW0Xvd5n+KJOrMeTu5nkF50yF1Ms4nOoajH8+
OOoV46OtaRmCHUJ6s96gFHs8/Z1vDI8CHAzhr2s+rCjsTIwMWyimHWk12pjDrEEASOhnhi5Nv6mq
19WEHWm5BfSUSSq++P3tt2NWxlMcSQoBjffh2t5iH60CTTQATxF+jujmzmCEjgKCL7W0DLWfgoQS
RpK74asj000xwMqCMx4hym5VsGgL8ydiIh9hFtsjeEle+ePXy5tT+bEYxMK8QjgvYslgqtkEHE1+
isAItd0ToAunPAkd0uGYSFbAi/Fg/piXVM82N+M54LJWCZouX6y/cjK79NUIW1p8dZyGpe9Piqux
9RF5mjzTmNEcJajTV2SZ9LHy3rt4yrc55dKzOVoLVpCCQaGWUpfAm5a6XNWLyvB7WuzGJO4xz8cZ
+7Oy/kXbtikrFovIhyeQWgiU4ibCIixIuylzgVjaPfrHp6Z7M5O+thLkvjtK4a780g79XwZ3aRhD
Ck1tNNExF1k8C7F++HEBPqAl2M+hj5/RZaeGgxEeo33MOwEiVQXBTQWCJ9BXwOTrqWXwjnQ7HkeA
AgvNoA7JxBY2W+LuXwePRMD8m42fZRy102CRpbo87YWM+CXdyElQ2gz2hNPzuvxZh4NRVSMsUcnN
KiHUrRaCVJtlg0Ad0KX78zvRW5uGIZYBxYHW4dsg7xMo0ckAjOWw1YZvibouUsB0C2RYPULjMXV8
kTVlhPxqZEzr6VXQjx2o7W/vgFLslZoUbNrdF/+R8CsRk56IjWccXQA/kIFulczVQgC8lEHtRaUH
+kz9aZEgARlsA7Et3aIeSxDZjHB+IZQLamx2kpwMyHtkrmmSW8HhrC9l4/q1z7Znj/balcrecaWI
oxbzs2+DAyGIq9321Mgk8wGwfJzLQ4EyEKVjVqHKaxacYw9U/KgtcYYzrbSSczfE8CX/wQI/T/LL
GhTP4PQrjQFbb0WSei2BuA4zTiYCBICq+tAsPBE+R2BLo4O9XIKpe9Y7xXc+x3GUQvKDbdIYopne
0M0aRzo7+UBa9e5LgFVgJyYqAWl8fgedYkzaxUh1Auf7exmedETFYTYv1qzZ3JaJ5IkQf49RVX3p
f1Zv1qBLi6QZeiaMGfbVB+sB/lTClJBPJlz4xHCu1KqUoilvh49PL+8HpYGdNkyPi5xc9aV56M+B
Uk3dMu3SuWG3YhY1yst0GPmpnBq610eBOVTmtjq4KSvvHs8RVb0AsBgMizte/sqQY+p7tlqmbBWU
SicGjUg0Oi2ARnyWKKzCkF0XwJQGuMbQ2J1/ZQk6V/q6eZo59jTDSBFH9jikE8J1hxWYbkH28Yjf
K8VJ4rNYacpn4exRprfm8BpDi7gsKyJLFe3JWlxTDVeror5cAvrjU/zWBC8tx1y1a33K5X093tpO
EbouRtAOfvvbtxSGkfdezNl/RDn2WUVo38kzikfKxpfBIAIWfehfK5ITBpIzODoW7Wkimvvp2a3S
GlilF9mweuP+oMzSV20wzc0E7mqPAWVvzD+VeYFMRNKX4VzsK/vE4+g5Q4KJI8aupVkhjXBtJ6nP
DcZk535J/axhntViHnUEn5lNRLwtVYYVCms+jFKxtbzT3nb2Pstbw8QSBoFeeclRdztIj8OQtlyG
ehLxWklbyLDCAnWHOSAekS6P2V5R1wbhbRaDu3BXGjtoeen3Mm5HCWI6bTDZrNucO71bAJI+W7Hk
5YIyYX06gHnIWbbsopRD2kQ1OPtHEsOlMPQZSSVrCAfqAHAIsfS/QXwowdsayTAY5/EBJRWadNdC
JAsOwAb/LgKeM5ITm0ALxl6HqSRXi8iMPHcuhJ/89eF4tv7lGio6kb7vKamiWKZN0wvU4w2lOUK3
rac7KDlEFuy8oHH/7RX6GNOzJzrscnI96d90ZdvnUgOm4Qow4EIuATb97PDVhMkGfJIh2bdedLJa
0/TJSFbi13gUz87L1TMFJsxvypa9zlXeKCMjoaphmOsmHyOwSbgL57TbYt+XYRJa8iMJg0FlViC8
cRR/bSr3gVTe9mndRSkhDsYL2mRTL6RdkePRXZVmPWWvgfmal9CoMBcluo/4bqqDFlpCjItx6uFM
f6y0mqirqa/Zms0xFhGcYIAQKprAl4Q4bZ4Gnnly78hagDcqaU+O6uBRfuYLySY5578zT3L4rmHe
1lM3F7Nnnb9X+gwjyqtLDaq1prQ2cU9tSnZLf6owl893Pv4KCKcvQOJQXRKOV+cp3vA0k375mL0/
ul/WmmzQo3DfpTbEyXBM+V19hayLV5rbAIidv4nP1NuhPffLVAO9EXE1mKdDj64GZD3MoYYbVBVW
oKc5qEvHh0rChQzd4bdOqCVNY5PmRtz64v6LQhmw+c3QELs0X2yppjIBFbtv0Gh4XSx0aHNV5u6M
TS+9zFR0iTliteDkHveUfCleXQnW3rZ0y7E85To9eXO3UJ2JmgFXQJnTAWbeO2Oso5cbfuukcp60
Y1VgjQqAoKQ0uMDKmMqATS50Ar/3Gy1WjcdmkHxOmcuZo0GVbZVSHIXBXTqauv5J4sShonZsra0Q
PsnFekJrhH0Ymg8FMhB0gHpTCaaOa7KcbzdwBOCx+WJn11kSjbxV9bQb1wc5S5XeVXA+gLqy6y4g
HNPfrwTcIiSjiy0xX/lztyd3P5iWC5IeY26tI6f1salZeISeDufU2SNZIdLwqfKhWvAIKyZJ875u
5pcAuhP/1wJS40BpC36XCmirJI2DieuBfXrzTWY92r+R9KDUYb8BVrFYkaHFinvzNyE2G9JZU/b7
Pw6PqhYjWyKD7CwNHO0hXC861bme0cYNkHYFqimHZcOi2Jl6vsubgIPaYDaOHaR5vvW9bdg8b0ZA
GpPZXwtccYSJ1erHDBf5b1mgVLvbf0YvVWi3F91LSLW+m7Ma1g2T5jiHXrzu0u1ZnhSswFpiLStj
LOai3pGGzg4lTHuqqzMI7FSpQ4KMFCdCeI5aYEt5qyYEC6HFPGQeIGBsd1DA4zWR+Wybj6GFsgO6
gHfOKR4DwFgjFWmEyZ/7stVmiJTxPwOpdRN7wpZni1Fn8eJ1Jrb7VlObSFb8s+z1SmgzQIGA7HvR
ci5OrykzFKoRYi/4wPg42X38+JQ9zsqvGmDWRkvwc0q3O377X+34I92OchIACcXs5sS960qLfAES
BThasgbpGsc8BFIidv3q7LTOJ+1XZaeXPUSiKY0dkGCc/8hOZSzTmR5wYyu6kj0QqQ1oYTKf0AWT
NsGsjkI09o2lnvc9Dvrzrg2u1j5FFPcSrvP9GygRhfx9wXmXrEhlI9IBe8MjjrVcCKe0qBB6UDgE
hRWk9/eQih3Vt48DIeRPYQAT8IDcvtVvtS0ODI2C3xe5HNHqf3q3dGFROaczNMe66N7BeN3GXxks
TiNGdamyZNTa19GLm4sIrnsRamDcUTPVahKgy8gNZ9OkT38l+YIn+1pX2C7k+ALmJmUEPQaI57MO
iD9dPncPgSoguQTPtWwAapfZhQ774b7T/6wR5f9HCQS3igIyKwLwT+EOoyHDlFZxVzXWMsBI8RPG
mnlCBArOYa/QCZmKigvEsTkb/90EtM0KF+GBxujcGhbNaW9kNdTu3/VHoHCHRi7CD5tfgW0m26cW
4oD4ObP+C0mizPh83f+VfrBk7KwCRaOEVKeRyzfAYuVJq7tQ0TqI7yqGuXoBGSaMnT1xeVnhT1do
k2miPws586pzsmFe+gYQoHDE9RnK0M7oaQU/av7Ebrjo8L7FSjOk/Wzj4WlItZRJ/vcSNZMTzK9A
tzbRiJ/SCCt8Vk5QCaSl6xffj5FB+loeMFljGoQhsoJOlb34n1wlSvFpV83X+tFmOC95YDnL6iMT
yd7ElMS3O65UZswLF26NmJt7J+Fmx5shocaAJWoO61bFkOJF2IgASKbwxyY8f3jxq1wAw6tTPe9p
rHgRSEzNxSbtD+0gDTRG0KQjngiCJjoQgrfX02Zgb5OfebBGO3T/3y5hvNGREVtRn9wg/KPrkY3t
Z4xlucNg56dShj2whlD4YvjNq88mKKV9nLhFFpSrH9fE5mqOZjC/YoIEQ0e42lMWoDsRjLRVlXUD
CnphJSv0+5gZx1AsOvZsCk1yVHe0UlnDIUEHPnj1Mxu6uAIvsvGMp/8mq5h6gDA01VFQuFwe5wyO
bLrpBN98f0uE93750LdQieN4WDoUikYZaIyME0B9tAjLpAUwHaC0FwHuFpEVjcs58/usLOfAcCeo
KbB09ht8Uv2I9qSBW4c1yAacomTmLRDZ/C+DrvupcaD15moc67pLxYV/+7l+RLvSAKQyCOXiSY+h
yTfS04u1kPaZ7kvu2+pZ8UeCFSeFPN1DPhYlHnm9SOmIxYb8bR3xNNS6cUnf3pMrOWtLdMaqflJg
+yWSsFMcE5KSP5hvK3HdxyPawZ+kQ5yeZ6D7uHUEt3Z/eG+7WbN8k0hImPI/PGI1tjM/BQE/K9qo
LdN+aW/N/x7AWGlkVndjaL3A5tPqDy2+v3OVp7nc9ih7jS0rBNtoSQkA2B0nvIq30egV1ubb/lJC
/KwaevBfpOYJmhVICXmZV20dPYRxCVKE8EgSSLlFnqJHhL3Wy16xKhVYz4YSePY0OuTTE0aEZ+BC
hJxBj6NGW02vkn+k2UGrSFSDFrXsPPINmhb+0RBQwXEqzHvHR0Q0JB7/XZxg1H/iUSPfO5NdHP/F
nJ6W+5tX+FBZdlUsqcg5H64ZcJQe2vwt66Edoaof5sVjxyTvV2xF71xjY2TFINh8s7qIat+3ksj2
mZTRMVLiXbKFK2LHqLqb4uC1LaqRHZ9xoYNeRBkThbfmQO2blOZkjfDd6osWcrUpLY/woxmSqpPM
OK1u17IUQVpZunq0KRF5GswC+wmU+hxRAoJsknv3Ju6aRdcdklU+WN9EmD+oLZZL8yuw6MLZHHML
9lO1XOzARitPQ9uVRiVswr1AGsf+kUBz6QPpXGtceU7vMjD1ZUCVTJ8j6LP3gD2lOTQY8WH2uSYB
5GYnq80PJJQyv4xiSdJQPe9wugD1FH0kkgTSZhosMIpXKU4qBNqFX+NWmogKHEF0L+ODop6F4ajH
wrUjo4dAZC6h+NuXG1AqlurHq1Z5L5NRQ365rTMm8bKMt8/jn25TlsoYNB80omB5aV3ar0Oqawm7
Efq/T2hOISqPBTvezn0vKaHuyL0eBBOnLYs0ZaIGfvL/ns6Occ68UZjEgpoWiXb3Or8URlmULdEf
XyNBw430tgoRNlocYxLIOHrc3Ijgamj3JPiw83Dm3SAO/DFN/iRZ6K/pEThQGJrBzypeDpKe60MB
eiK6upPtg/NEC7vj6tHvq7bbldO+afX0oHqiyjjxVN6HSlhZtp47QoswGfEulE7rGPClTdO1aJ5D
lvwwU3GXXKTfLqbQ4qHwSzOPr9WrFDO3jd7vuppjzjQCpkb8JlETzNlOXVfOcXYdWqbCIG3XCTpH
Sv7/SIbh1oCQjll5emMHsPQE8eCzhrdjUkGao6hs8tZMXnFZh/YuLIo2rJqZInmg39lbuyY50vq8
aYzQ/zWjcAQ6Mitvzcj8mbEYMFNw1Jj/DbieI7/aVCiUkCYeV5o26Xc73i5NYChUpQvLFhiysCao
mKWk+y4owh46DJr+ApijojnFFEGe9/wbNWDjUv/S8MhO2bq2u7LMCLzA4KMXqakmT+iZ39x94vka
1xdDq8vy4oS2OrLcSJOZ+vOjuN6zwlsQ7P2R6VFq0N04bLw38wJtR/AtTC2IsjfxUga3RQDurV5O
TQj17vQdLbwuh3HK1jSNmYpde0XZA5Rjs+H6nY9cg6gReFO8RuYcTUxYHTp6SIzmfSTMr1ytislX
hJCObSz/ZRpLWZK4PMhfhNdDArxQTtyR3YWTq47/4CcFVn3WaZMiDok1l1TiczWPIrT2SznKNdnx
DnkeN8ld5d62E/5N3rkiTmnLzZ3BWegmkxHAoCj3kkOlUy6Hg7A/U6sWkEP38v55tD23idYAFHz9
tced2OApK9y8S5QJOOyRCO8KpdHzAjKZAOxZRRxKI2kr4D54FlqYP8BECMzQWGuDPSgDIs5lOHKF
e+ePpB9wVoOAQSN0eHWgf7/tgM7GHmvkiUrwYDloAlYNL66vWgJJ2SEY6RaD/FF3jMLYm2LpOW6J
P6FPF6723rJ/I4VGHQmGfBWzRJkLJ/2goQEoGp4tmQbPzorNQJSBxmG1jKNznPzJXQoL9TNBoDUl
MI83DdmLpS2QAtzBjwUAVBJJEDxq/chYpR0B1vDnTIrlInib8PFDkIIXkacBT8515OWrhRD2QT+X
BtUIyuhIqEWAwUqSsmBRqSW0LBqBShp12Tu++K8GHMfHUWZNyoWS7eivPqM5YPdcT5vVVy5PMURi
h88QnwOqL0kZvKiW2Vf43tI7ieY5QRq9r2RTo3+cfzPl0XFM3aJ8oHLy04K8ZI63CtTLGho9hbnf
avXYf6ssbOLa17EjlviVFvBbtKx9MRU2AntqwiuaJlI3/HDEkI6vps/tDlHE/FV8AaRRrP7J93Qy
bHfWwn1jcXcT6Uq4oDDMOsIZOALumiJ2+O67kSrV3XY0uP86tEpgSUmsPPjO76pfcz7d8jvuAk2T
u1ZW8DJezGB96XFE0sVDw0rcQINMiMh+wxCWdyXHcgQXVA6ctdBCK88CSJMyD9IGg+Y1FUDQ0XA7
sN9y0XrmorSd7u/iUaop1g9uax6pCOH4XRDhGMtCVSlC42Cazt9XHgVV6xGXXZag4TGAI5y6DYTc
h2AyaOd4+fqw6r+sUsqG8fQHK2oXnMgAl6nzDAZ6rDaPtuX2y93ryPq4VzEor3ZVOHHYdmGkyPb/
UjdcnHWiORtTcbgPm5zM6XYKgEjYvpAxLe9Kvt2Byh8pyr1SIzxbQ/u7TNRSCc0uloFkIB9jN3gz
qRcD5pGql21Jxgxo94BvlzJN4p1Hw3NodbtxTr8B3Kx6hXosVCtHJKeifqAQxr+MpQBpYAy4A5TJ
c8kFc6igaVZsT1v9UQOr2Z/2DmItNniBK7gfQ0MBPfInz2SdgO5dhTQtEXTwiYfxgl9MfUMORB20
/oexg7Hxli9S11bn/8W3r6f7licBTqOsB8X8XxMOu25+eI0YawuEmEKDibf4eHT6B+/PdcsuyQEV
K2EnQhQCMirrlG8h/S+07YAT2OvqrsumecC7VsINpAjJ3gmR4+32/mkLaEVgD3rf5ZNGYwpUYU6K
gYFdHj0rJ65U7PU7pNPzXNy7JzeghL6T3GaCQvsQ8umzw6lcIsHyhDD/wGfS+U6yRQvL7Tfqw/va
ojrILb7y5gwis0TndT062f8N9B2Ot3hqdd5VOl+cznn/fh9aELV/xwRftwgcYUbb8hoasLOw30Re
4Kq7dGOqGMCm4fR6+Sg7pYs7U5P5E8HSB2vUdq+dQMG+adANS7d0fGr9ryioK9vYD0MVBhJVrCb0
zPz9WZdeAxuhJHSj6YbcuK0AtKDafuI9V9VtEkjQ3tjHEz6zlCQKwlAFtdRBJe01COYwoU8xW1pt
W1tVouiB0fburNRjm0gI8N75WJKrmEwqgiLr3m/Yrpp70p+8NDnhtNxc3I/Nby9lpLyOxsaLIuww
rrXXWiale6uOIa4VKzIFV+6dM8qGj6yDdP3Ym508R5Ig6rkV5BzOc6NtkxGPGW1PV6/8ZlaV7y3A
3yT6E3BI/7IVY2WHiFpzIfrmgX3lWpcS5fSPabTE9YW+Q9+jSRg1DJ/+Ra+FScfJBMJTJo9O6a2a
hTza017aIsAxDakz3wwYBazLnC8UI9vBIIe363KReX4FVyrLA84hqAT/j5/uAh3Rk+yjIzmgx0GE
nRMvAzYfLSaMKWHWkzPFqSX2L4rKzNjQbiWgglv/RSophMYpwozzoU3yGImY4sWhC0BzEBYedoWW
YNVHNqcFSAwqBptz3CXuAotUKHAuTsNWno6XnnpBTDOT+Z2UhhmnkGjDnG+P1D9zFcd3y8ygXfI6
HwJygNCJSg1xbH/aPOHG43dJl0myQYTC5cYK34XiMNjgkAw/aedTR87caiF+V2uyEfINjOm9a9iM
/RQ/PJF0vHQEsEA5r5ZwKahQb0cTln6Ln1e/p/ViY9fFjVP1E/ANmA93xtSjfaycm7FtogBn0V5Y
Y3y/jLoLWqC86Tk8zia6OGxG5R7xqZ10QPevrK2esXYOIxepoZsFwi73UmqJ89e0EE0bp1uNnvbO
9TEgMNzvkuxiqaMatL9xFWCTGwpYTunWztBehC8iFnDXtVxhHxCtCsVtWPYR+olHyjo7uz8IS31N
T77HPMJERAGx0f+idRQE7J6VvOv4ly7OyR6J3RHAvX6C9WpKMdRzG0Vlew6K9ZcN2ogzersdpwRL
athy+YwLYji5HA0mb5wV2NiS93jXXw3v6Sbx5YPR8a6IDA48fMppAa2yoLe+Ai74puRZLsTuolEj
9/iqUC8c7dw4Lm10d3oVrbTxOfExV86G3jqNzUK/EeY962niR/dSlQ0HMa8/+6WZg+NZbF4fAAqa
/LCKETkSepJE98UjL5NJYNuMNAUG+8c0eAmWvBIkCy2uTk+CVVubCLMf6Mj4si/UJejcLH0UsPAV
AKOfQ2lFoPU2Tu5zuHz71GAx0jest2R6bBsCcT/+26nJGvv7i83i6GQYovXSoqHLDH3H95IqYJeF
HJz0FDfWCbXOCbExXpAWWHFEJIa308edzVh/TiXcjXtu4MxkhSpitgFLm6vYE53Vlrr4N27cGUvt
TF/b4Ei/cBKsua7F7Vo4tsAGl9/rIIcqNwA51VaOOTXTs1PoBZYiegs14P0nlNSenb9AtKDEjbou
iYUGECiS5H+mY4KOdYnjqQ9UmiiWLKjszI7EwA9C6mtVtYtUdUHSVMTSDrO9O47SmVl4Jp9R4C4g
Q8cFBDCFnmNYiEJE8wFGMeI1Gjf0OgqSjKJgKhjvGtnzgf0t/+/4fObkjm0gPjbT4riyXTTWutOm
qCVQrHU0coqnGnXG68ouG1fU5f/5BGgDSg9vabNXVh5e/4X4hYZSThddSBusP/0gD7TUNcXOSMyc
m/Yc2prePOjZS+KY2TyBKLjNlx55ZD3D/T3tTUSsps6YS7dHWd5Gz8yifTIeABYgicOFATTy9g/D
HJaEV5aasq1RmJIKdu586GTCYmjNpNBjbUzMhuufVZ2GhAOqsOj+Co1pFqUX1y7STIhCmekNvOjK
bcGF/jyEh2qEGL6wbo8qWjs9RK07YCDbtlq1CCyXwz8+VbBmbz2JGsuHHAh28JtbWpV7vArGG4Fw
FjesfxRtkrWvXbnoz0tZ1HAZX6BejfnaPyZu/Yb8UoG7xlJnqkp2N+/52hvigj8daTAUaYD94o80
ZZkB8qnpdoGQzwBbfrXM6RBXkbODq1SYYKZ63N5YthbgqEUzu2sd7BRIh8NCEvcF1uoAnlK8lFgL
pukz9dgaiYwdsWwEhzyUIW5IxJer+yhU9iHCcWLCBLjLOH15GJ9sdOt/es2oKwkI1+liu9A9wmdU
1TYErXQDP27DetyA1muzLSU4leJ2BcGez6l9Hi6Pk83TAxTDJhSTjyloW7NM4vLCqkZTuKCJlR4t
UAp7E4/UtO2O2eC2XgxQ6AZ8ioCUgjTK65e/Q2MO0AYqWA/1w31uDnPYDrnRou/KuECnPxVCEr/r
Ie7OEC81QmGYmhVTPjO9daEIcl7j8c9M9Q8e2zbsJkQDtgaK0bjLPQStogAEGLedbd0gD2p008hE
E/scycHNiS7XMk+MMlT5zOawZrLYbZOLH29Y9lb5a+AcD28+lN99y0zH3li+RbOtfKfzOxa/irKK
NE3i3jCBwnqRLweBBDFDTQHC3jGDtm/A20XRyuln4wtS2xsOXvOh/RjtcOlOan8nfVVWu6o4RJPb
moogixaOy69UDWgPgz3EBy/uov8lh3y5YaevszWbjOn/wedXgVNDDiAS69IVaqFkaM1+O3YgDYt/
/mZMCPOmsdbmRobm2RecBFREPKY5e8L86iR1a9Qybci/MMnKCPCaaY+OUc8uVmw/WgIjlQjgxBch
4VW/8lU+ay72VqoLT/sDLrQ4G2vYuJqS5GS9Jg5+gSxtilKA/WneTiUYrmGcf4E/TLobxNYoge7J
lYyGTofRcVTjLpKut9XUoW50Hvw/PcQHM9Gi7Vw1eiocoQfWiJ7mg3yJ09KzzKYnU63c01BaZijc
5poCBAgu9pjZNvSkJQmiXb36ClOmvMOVZvzN4L+us7zEfoUdI8Kfhj/E+XScqZbonn/Ye4P10Y7o
vhaRUMBd5xhQQU1yRHaywKbztLS2JWjJqrtpEcxNsMWwIAOfbWAV1Hqk/er4ucMtujndOIhAT4OI
NItMv2Uq8uJ8WKyMDQtOvNnkHKngGZ4qDPVBAzzY27aRB6pznmL1x+HgS/6Mk9uipcuPsUXTARRB
FR0F1kF25utdVLAJlO+TIHWpdUE7dl+uN++eVTEoa1u5Fol9ugRSXOwrKJpEEr10MDX3gXIGozmM
UV/ZAm4r1iOrNrinTJum/nrof7JCkjlZOO84UdRx1XKtlCSZc57HbyZ+s9qOytLqb8C5riMTjFK7
mdDG6Jyu6+a7A5qAuG2Y+LBYPzdTIo3gIZXVab9HChB8TuPzmlyg/QdshbbkEKDJ2D0sn2IWvMIZ
gwNrjYLEhY/ADBIHg+4mEJykt9s9JkUm5pHJLdDfc7/iJUV7gMMPp4kLYpuxZZOuvGLi/tNgcFpb
7bjuWD0g7CyvNfZgv+fYskOC8VC2lwlOMN/qCdFz/SUg/By914cCv8ZM2J0EUUaIuyDW3cIHM9Aa
VfHADGbSEWW7cGQtp+px1QjKysoIaxC60mP6vwHQgkdaUtU+Uw8g4iGNnyswJEE6CKptn9pG3Fk2
cD9Q4cXKedBJ7aZbbBtrrJMxuTzJ6bxZ8DiHDlbe7RNVD8oQLmeugSEO9iEyZx58AFv2B88FP7ln
seFIxo1N6g0CZASQwXxsX2woyxJyChjXY0laQD8JVsDwB+K6YW59y9wB7AhmeUikv0vsnSHHKwYn
m22oS7rYOORH9PNh1f39A2hLb4JqfkUT9FXIp7WiH1rTKvJLmLngUTfn7PnQQOp7aPeFBWIsehfD
FX/pLJSK/pdkXGFzPd9affYtzJ23MENe6Z4mcQaHFN7MkMZGmaZlRwpICgZx7XkcJLbSRWa1YqT/
9dkARhNQv75pauvVh9p8TndBoOW9QYZeXqG5iH/u6Snp+z3kcdyZCZ/Bejq5wy8qbNGSFP65LM/7
84Lp1L9GNp7Yx2GiafspYyCkplsHihsOy81HSzYVXv26STJ9QHPgKFUKHDdg3qKdJhlE0jlViuM/
Qv7ni0gG5CnYe4yWFPvW0GCbbqhX3ZkhfhdYrY/TdImRcivzAtVPdbQtqVeGE9ISD8GqpVqP5QoB
RI/bdGbmLMt0AwDOmoFR785+vcg1w505TP92hdUrVtNq90syk/RX8KbmruD96GjbCk6isjWogjyV
qK0KVkIFSu09F2XcUTal3Yqr08mAIEsefMSVXMUdPFUJwYIpr5t6XhBrH0HQmWfFGWf+30L6BRTQ
Fa1B2GnVqaLbAM3vnUXUVrv+PQkNsgtxlfXnAPAUQNm5JJf6BZt4WXDfuzS4oGhNRjGXaz1qds38
oZNz+bOHKKeE42XJ2inaksu3MTI1QdW3kZk8ZnbWAsucvisnj8F9y8L4c5gm/M2hVes79+bq/Ywz
m89FiKLLoMwcaNSFNryvVxIoKifu2YnLm5Py966XSZ/zV2LxVB3+tldKUOZvEs2+2Nk5oLwi/oyp
9HV786WER3IyxbxqV/bMMOdTHvmURCFSBdlirMSbwwiFWzBrSJ5CRORr6IBENlxf2TFhl9n+59/Q
5ZQWsZzDLpD4758rxidu/oTiWvjuB3JfwgZflAR1PART01kS/tPIJyok/NSIrT6YTpDbiXMdKFe+
xTraZOaRzB1DQv0PtRr9krJL7kX8/2T1Z/OI75cmzThlVBqW7IoaEpz9AeDw8QDGEet8r+6F6IYx
pXMCFVzR10BnlUltrzx77IrmWegeHcnJ/g32NgkksxyN6NgZplArGR5AVwYWpLjEQhYATdHVjT0E
XC3ant1zsyLOYmIeN69/cF5KKX0o3rnYGDrpkRjKgCwqA+vcs2KMdF/zYwclxsKZWF9y2AK6gB35
sP+RlJjRAR/v7fggc2kYkBvXAgnw5P1unUAu2x7Q0tnH6iIuTZz0Bf5/m4dU8f2dsHrcx0Qc28yK
0IAdcvHBJLwdPLOsCb8HH4gdP1VS033UOlVZSNoPN65lYhXD1V2LRg5s0jXK5QeMOc9jdDL+sLXq
jJmFz+rngyeF4dWfcSf2C/akdQNRcq+67CBHZL3HmRTlSLd/giJ4oISIPzACv7jVqSsoR3FiOA/P
OPQD+CBa46156VGcLcKw+WMI5JBM0nogSwUNVdBFGu364Eh6bdrN626ku9erZ8IgJ/ZFtjViSYFg
vxCZuQibVQFUfBn1xEzu52D7xiJOt+U+BNAEoB780j+DAkgGJN4XcBi4MqSf011I+/hv3qPqhThx
do0EzETwxkMbYh9UapcrZwIV4I5FnPoisTd/GeK2lih76+qlGFnT/YaFMYlzu18mJ+301NV9N4/y
6kOnT5e7l9q8e2kdmZYCxXFxWdMMKqfNUo1jU+8SADtRASpGHaNuRTwZpQjvR5kbd1toYeGmD/Fa
nd/6SIjdlWq5W4HryZ9uwzPx8XbIPmXxGpXj91uutotdI708i2fumiPz3xTMsFFqnMRElUiYLoEv
2naIAgalXSWbVc/N8rYBLiOF3y40m2z5duuRsvzG/CptqpI5aZNVRSjAyveAX+ojBFnq9Vm8hyrw
7Klu6H8WPkkmhic0I8GKkOejZOTbfnR6CO+erN8JyfvRVUnen+M3RCBteVklSe9572ApEdcGcDza
y8pCxHeJAB9fokiixraQF1noO4SpIp5skTTzcCOqL4ylqy8oy+FkSwOr7dyfEen6b8sMU111jPwn
elEE+SiA7XEW05p5Ub8KFtQbQO4BxIj5XyGWtbvwgL7qnLeGWTj/KjenY/DdgqkEApJ1dti5fOY4
8nJOIiLGEP+Whqu5tYA2i52Bv93fI8gd27SuorlDswcwX/5mmVy6h6s1niPXauW3b5NWsXM0mh/v
3GQ5kDKg42wxPg400AqX4aaM0QvgiqCUx/71RREGRooChFvhhiJMaUF+96hUUSAPqZnOxDVfilKn
OaL+x0EQpIHJZnaHD9lix37LB2XaXdL8gX/G43wKOzEmkgxJjyfRm9iui7AX615NpOGLh1Jdc/7P
y7Gn7JwpL6iBb0belydEqCjFyJ5uqWwOFqea0lUaOdtNb3gyRJdhXM6Tcwlxa8Sq7w/qhuBch2Vl
ueRbWMIZE5Cl9tVm/adQY68gHiQqqYdPqx8jRvCCtVtTUxPWQOOn6+SHdax0IL+Ku+F8jsNcytne
pKNrxDCGsmBDOM+97dV6lM+8byPozDKFnhEHee0fn0pNSpsxAU3j5E8T6aK1OEGYgeenGCtpVXSX
/uqydgR26VnOMCWXyJ7Sd19A7xUXK3sGsMpNTsJ39XHCD1R1L0tw1SG6onhVpoHFGYbMoo0Uhc66
v0ZCAyi6x9sk3giRMUElLo1vh3sfdeJnLHz9uPs2ZKR/cWkOudhP4oK1q9diHQS1YVII8RRJ4zWN
JFzvs49ucPk48Yb4ZCEIzD8StOr3NHEIUQWbOWVk6zefl8ylSyOFTfl70YzkCwPLUQg7Y8pqidgn
scaZIL7TUcjRzXP1/vtz+04MmwN509GkHq3iqKmNt0eQQID1xNqL/e749Hs9nYIaZkvSMMBIcRAP
SKB1dz+iBys3xHzbSNUAvFXntaT6bd/i+gI0LA4PZ9yOrkpxrGndt5/CgCgUZUaheZiRmXq+wMoo
EtYvEdV3tug5rP5q7okZJZh94wFHMUXVZi2qsjHRENGKurg0WbBJgQ3Cjxd8P7f2ptmFw+FpkbIs
0/ET+/Ac/Mb1j68xkLwPTPTcQmVetuEVoRu2yQGicQOv48DK6OC00Zr69Zr+3zKuKsoRtxp30iIQ
vjd+vrxwmCQgTvRTUEkz2vWiyjXEJX3Z5qpxxPM/OkHkGmaxLgGzNOrB0fDE4Yi3CTawjje8RV0v
HISqVyo0wH5QOcZWlPn6/kAuYAq9/UyurRmUoiR0sb5k7FGF2rHjiHhVI55C1H3zovzlfVl2RLS1
LH/5CaEsd8Qx6ATZaYYLd15OxfjU0sEZXZkbuAdBDHZABpx2H3EjyfA6zJXxYSe8xhtzI3KuF+4X
oRt1dwwEiGqD1bTHgbLkyUyda2AXzWIqcz1JojFRd9Z1mPwSw+TSjO/C+urssjl27hWLxg5stzss
D9mN1eSdSA+o5f9J8e/o4PPE2cSs6Hvh/ucJcgJGD7e5AAUccx2NxsDMgUwdhUdRfu4DYv1q/H24
vAiTX6V5Q3eDgfL+LBuG7tv8gNxLmUQfapaT0yDvP5LXvb0ehtlp7eqyBAT7o82acFegixmBljhG
mXT4ERqVEkmsgAgRPs0pnxjoPg/tuRsW/0gXe/I8MVRlk+IIBClNz1Ns4nUNG9CMpeehZc1SJDSK
r/YK+YuV0EPOzI0fgjQxQWi46HncACDdYcwv8fPwt4/ffsp5/ybX/sj3DSqmNDFdQGd+wRKB6LzY
EvNYdqBFSbFy3siCH1vbMuixZnNVbBbekPrvx7FQiHzOCOFb92rzNKDG7qdCMCAxWUAjVIsVkP7n
wNO23SXPGMZptMr/aNDhF2vt6HoqwwZ2GPUK/GK0Hn769TzWvfItTrLPFYy6QJYXogKWIjU7j6Cu
zOzRarJ187FaSPXGwRtMuQFBih2ijQ/JRRN9ZsJC306ufOmI+Jlvp7NO0PE/tz5cHBdjQf0EZ8k9
auf5uOCedRqJukfAcMS7TkGbmynmFiVq9HeLIPTqtRgPE01FrJ/7Tr04TyrVKsSSXQPrWOeApDr5
Y6GG6TuKGRSIN1alSRLOU+BclNjSEAW1deT5mlTzg+Cqcy7ygM65xoTCMrLteh8BHD43qanyG9O1
7JOc0C5eowuDfJ3U1c+dAztphdr4bkBAhrIPzXOQqVa9IAniyYP3HaCvHdsFA+rbg10rUs4rlBsD
9SQzmrJC2tLIlfUUrKSswxZYDnYaDbx5QyO5IO6jHVKg00/9RCghwTt6BYLC677GyXp8yi7w+Zfe
J0U4UGGTIq7FZzE9TlFRypmc5IXVaYX/idRpiPGCylVR5ppjHg70g8q8B4PK0J2/tr89R7RM86KF
PMpBG3WyVkPsxns3d0QkfW8iH1kVZ1xkfJg5qfBvPJ67o+WrboOY8GTA9M659WSDUEVeaJsw3Ehz
e2/tiCeYcvHZBPXF6f7Q6FDERT17LvxFYdOM4Mrd3jIuWniGLbb+TQm0XoyYjSqQlb7F1xtlpMqZ
0NeGc6tWoqB9O5FMhR6p/f+NV/9bvVgtOljIcxiFmqfT/XfIK81tw9x+2jJq8EIV7KRtuJa3T7bJ
lVoV1VubSptwm619kOg4Dds5hElVAErAJvMXJfvZfc/MukLqOiEBAvzUULIXRb/u1M6mUIWp04BE
8iNqm8FDwb9qIsR+kfIzAqyIvqvu2WR9RJ66+yh0ByEisBILQYduoVXzusBAQGk4o+ARaikkBtLd
oS7SO8b1wb/PTBF7QDs6oA/nCk2Y80EB7EV/VElBFpc7Gwo5VJ2wAfDuI2/iWSQVM35dSFN1to4N
aADMjtg9gI4awEsTfApRWddUhM/2BzOE5Hn96P24nBr9ri4hiWCQlq7y7wwiL1uvWN5szZc12akn
SiqghRf4dSbFyv3WJg2ETe7DXR3/FtFiwLMGU/aYv+6winUtvPQTrAekpHQ9dVfw1M4UmBxnYVU6
p2hnRgC7iODlPMsJVlXOW26mBYcZCSxH1q0VVDV5BEIrZUb1uSuxq7ef5PLVTfoxIcY3DpQPmikz
YKBO3VoXyusckU33sS8Oc6KYvHx4UaCe0jXpU7xDT/g7hkq/HSKrFwpGWoiiR/wYh9t1JJI4aL8j
V3BMPuhRpJ4jgd+dJHgISz7HrswmfjEvud47dWxEvvo8dqQAUYhZM8oJNeP+X+isw98dNXTZmukf
hcFJHnelpwb6F67ba85LtggzU7LZeFxGcmmE9ZmwO5eLc/MkZg6etYnLVSBb01ll0ncflRt3CORl
OExJsFin8oSql2hF3rf+6t2v6Clro9sGGNW2wz6/mOTJq98rC+ODx/BahwGSJYZWefxIbHxaIync
9Rf94uEsqTtyEdnVIGHPvVw+5NYxb2VjnYI6A43xcEmNczcFjOGPHAuHUocwgJSGLierMs4ICsVW
q0wwhbgM2Pe0y545qIS+L9e+1pfCb89Edoj/yUafC1npiUIS25Ar7tyqI2+W6OEttnsWLIhtILpg
3k3+J6L7TlgNStVmltdB+/5nYJS0lkoqIuTm1CoIx4RbjsmaPN4dh8nM1kysMYocdtGdbA6zFJSy
8n/z5rcWuMVdPKIgxzOdTz+870rsrpztDioz8d76ThqqR2V9SzWUfeYBzZkt2GH27KidJrKhl9rA
EyaMwc38m1HhIPyJAgH/5CxTcC0U9L4FMVWCcSUZM56OanaIcFMvjE+iFGncoCntq9x6CSBII6ni
p8DR3IYkjzUY58q4J/MyyPBqV0FR1yDLub7pEfTg3I3bWLnbwf0z66jE71bUO6EXWHnPt8ciGYNk
7NmlUkGpPTvlt9++TXjR8MKTFgO0FTK+TVhH+tPRBBKWrzVHZWWXeCUOE+PhlpK5ox/JmblE4IrV
Yr488gkFpB/HpYPDboB5xaiBrWMU2yswHX7h7yXoV904cDefCVfDBXiHmwg1AYngF3FCqJZoJ+BS
STCqQ0epRB8Z6/sYN2jn3apfODsE0/sN+mlC8qY2lvAJUO6PyHHcKuHzw9SstbtWzOo3g4Hn/BI/
rjlFru5C3qkOOrx9vyN5bIAtwI320bHvNx89csqJhuilzOLwAkdEhzNMLkXelqrQ80w6H8iwU96X
vkOKnQ1IvP/IPh9uULH4R367Z4nH2vUCRoqLZio2WqJrQMlXtYDY4JNzYjl/RzNCO1wfyuSajwJ+
xcR9+ESV3vQecCQc22qcdr3XyqLNPHElYqMbNYkdkpZ7r1O0Kwke7NqWKRX5AZ3sXDyxJzY8C/nA
QBqjCPM1Yct0F9Am8uqAQBaL4eZS25t6LIYTO84XThj+y3ysXkqIi0NusQHO9SzpgfbOK5gos6LE
biwQjVk8unLQ5oFWXgQyt5Ep48HYrnUK1q6tMBooVWOftBNqZD85PBC/bMzekRKXMlu7vsLjHKtH
L+7ttwE9FHcJs1Oxe8daQKT6snVpsaCBxGeuE4U0ys0u23tRM/W4Z0gKyvscYPDqOTmIE007LR0F
kVGHbEyLwRlGJbQDFi8HQlgPKTAN2HdUWTER+u7vZgiIgg5tZpI/MI+bIH2iLBzXRVMFqU5iZfx+
L52T+4QdtUJh9VLvLGo7UMJMq17fMkSslYmlVWxVfeg9e8ktbX2ob/McRD4WgaJVryQcG2Ac1zmj
xM+20lV1RvIKk5BaLAu0zDTxJUEdXmACpg4xejTjDm2Y4Mq9tbc2qvQplhmiE8HFlaaT8dUHtWpP
z3wAD9tL3CDy9BYb4tfohoVxZof1oLMQn6eE3i/eJR8u7CZl09weOIPnWwFB87xHlY0KZp7W5XFF
bTncHYWgolimqH3bKa20VHjc1GJByCZUT+2d2scg6xZeCKbyY9INHDVLKNGr3xgxiKcsQtw2NvTK
yqEgST+ti/Vk4A7rwrbNYCTrKT9oKNxUVpL2kxWvEyevQeRbmRSxtuEnl//4O7A0/6sY8wLgm25p
PKyvVXBYo0N5RKEx9epfARLx6RZGuoFLrQTtp3B1ejvFB3UM6MXCMpznqs+QGV0K7X3X9wPOARlS
3koPKsve+ufqsRcpECZzUBcgP1BgLa52WIdtOM9dmn+JhLtHP2o82gOfHd1KK+0fkXucjzr3jRKJ
ULoqA7S8hdi2AUyk7qkXZsl+rAOw8c3rTH/9MxWMgM/Wub+fpPQpEidvdkvYytodKXnlCLl2mRWN
5A1lISjutWZ+y8QH2vQ4Rpktq5QsCKMQ5z3OstBvO228Nuw/tqt/9IoNh5VHE1NbH6DqztMYbGmF
orT6H9lcIGSfPoAXC2WL9rXk5eCmIyrEv1Nlyl4s0CBTdI0FdK8H83ADJsemIZp6beqL0DvBZZLz
XWVkzzbBlwUQrWR9qU5sXN4sjRqB0Q9ngmQAFSOe+q8WtcRYm+W7ppOuUgddnYO9HQFQgevmDfQS
5sYV3zQrFfP4KdeXc/ZNlvRFgwIQhWte5bag0+ehqxxvcDxp65pe9wRdQxDKOHbkuXHpmQzMHIiE
ybPIVPPGPEXV73FWxIDHMiRfmwhvQ+0r2g3O7jOJUal1Itt9bRx3ub4xbPNAVRNFJu/RZp68ntUa
QLU9Rx/bs4AVfznzJXKXq4L4YKT0RYJYTLWvZIt0u0EVhYvr35IqYmhzh6+3PZXok+oF0z5j65Ki
dQwaBAnQjVy6jXzzCCSxltutUBSj5TMC0E8ZnY3N4kH1qwluVslSZvNQ9SVJluBcsUn4LWnOcByn
XjfJXmB1I8/WFgNS0uiWvzw2cRmq7Ch0WyiLIXWruh/ZvNaeIwmbAaC1jMX/xZQDFFiaSHG+K6e6
ijtoeNwI76U/c4g8eRpKL5mlPg7Lb9hZo5Xbs+UgNFyL5w8wjEDYWYt0iDsZ5MJjyUsyN7JeVwZq
/xnaQidh/N8JMl77Gl0UkVh8rtS1z056xJ/BMuu1oQ/PsaKU2OQKbvM/zB0/58b6A9OyjmF/D/zC
oOsZVvbb18G3VpQ3Lk2JVJJVrwD1JYkcykxWyeRrKeEdTX9Qew34TiywxQadIkIsKvSrXam+akKs
R7wZ5SquXA7ErAzhlxivPgRTTnsjoVDjuMEytIocSsyMmWVtQootG/ISfMAa9fchKml7vo2Fl+dy
imuJruu7CPZCb9zmovCASnxrl3e8tU3BKrBTZdL/YFuFPsJpu5JLIzYwPwk8kDhfzVzXJ8hvZI+O
2ftBP17y+geppMfg705xpsl9fQDGsMSoFnZ04dYkMQQsFlQnsW9qMZpu45+NBS7x7tICdAtVGxRl
l6RWMosrHHw5eyF/ZDSCfhQecXrR1E50c5UTrVoUafClP5IOlbu0yjtUBONCfdButkXm0PvTvZ0C
NfPlCfi/q6RWzCnT19RyQvwXbqV7uDUa5SpJaKt/9iB3EO4ATq9bZEA1QdvwKB5Kea4dE1/i/5bY
sNk5K1fDXKTl91RwS09N1k3OcJHPQp4FhI9aW7FdEBKZdsA4ZUXwHQq3wrb8y0uhmBfcDTlBHY0n
IIw2yQV+VEXhoWLpwjkNc4Zfgy2kzo9PhDdT5eXO38J5lhveiRu64Id1Wixzev/2UU4qW9vPaimb
k+tGLp9K5I5465t0saaTjJCcKs5dq2nEMc/0TiYK3QSwQg0R1PAgsx0/gHaHSZHiHA2D/0+UwgB/
bfKC30M4Q7CHPfUPuLQH+Fy0MypJ1nPdlU1bTMMh0w7eIcI4kxzi8jWQL6llqpKfN0otmTVJ14Sd
PkpieAJOPUl73I+caaqc6yRq5J4QPO+pn2y5V+yS+hurZykgjxdMdHvFIsp2FOl26xsLMNyONTdd
bgWn5MEGndk3oYA8l7UyLFksXuq4fvWcGoTU5T/yD3wwnlqnc4HOuNd1RV2rVNDBN6+r/PBeZEMd
7ycxwsaobV3DV4+LoK4MvfFGREQGfa+b3zBmBGWTjNnTlStRsRWCDsZe6oJzYDptcLEU2TyJb4VX
Z3z/n5s3+fZbI1d7nQZoHEFsXhf92EMxjhpo4RYIjdr4MFIDR6+xYDA88GA4dsfarWpA09ARwM94
ej5soPXU1n8E4a1Xa661GFLSnV30lENf8TrcPfj89EhT5TxD4chQ2vCjJuessryyidAGBsxOPmBL
ttqfNnTXXGCgA+YyDIu817pxFSzce+AmW8eMdlD6yK5iQ/64bgQneawnPMzA8xwpHUaA6IIdjswY
x2c3dHot9GfDYPVp75J1Zq6NnWoQZ6xjUIMct9L2NiDVI8Vhh4qMpdN3XJ76DMCFJyjfZr37Vdc3
PjLWJ3CCnSAaJR7CamcQOx8eSVuSYHEVmC0gJve2zxvONy5iXyPYU8yH6IwyRwo9vgOtor/th1w/
jnCUl9LBdBywBWm3HKjtLgOGHx9iVxLNncuI7KWJPI5QGtFSVFETi2DMa7oKXXsrdPNC6S76gz9h
VcQgrOP7RHf7Hbsciyo52sBZ8/jBKkYfkTxrt7MR/jxCWlX83O5lpzvpC9x6C/GCuYpj1qPl7Rkz
aVcwy1OhSZ40sA8XeDbVTnVhybgT4u+vnP93ZeJa78/YVnMHTYNG1VRaPCy8wKRGhwzkfabHG4kt
makyRGM0MoBd47TqecitfiU+Sl/jBH2uz0Ekpa3LJK2LD416Aaa12P2qpQgSJUsh+rwwdUXwBj99
XpLabF9QxzNJ3/O8yUJ2Epdeab7JagpVvRn2xoHncUBRGsX/1OqsVp1qwHYHp7KmYC3fuU8TcASL
9i9LWrN8Dfz5dIS70Lw6JOl7NFaBL+sdcIbZvW6jeUI+ns/6PfisV/AXsGbB/5AAqXRLpdcF9IUU
9IIdBU2i2qkqpMaJ7sN0x6kX6I1BJ660hrbuyBRAWUPEJgUoVPhy++PpAlGlxEW8Xg8IzgANk8TK
CtNk8+9zM29wgcliLMIGE5BcqyJJsfzOLOffpvSZ9rBh2Ilg7r2gF/lFT0fT3OecM56mBnoR5HOh
oHgZXdT+i3EvBKkEyTxj26nrKVaTkYXnaV4CsWYljtosPlU0zaFKW3W4WuGdnGEQGEFS+VfiZHBR
8ijA+NHfXkcOyOgjlXhDS0VKBp4gsFZ9R8znxjHnJZLCP0O0pw8znUmed50R1RspqTP143857njC
mNbpy8T4U9PaaTcaw0tnACmXPpTk63Oczz2i+eQ67Px0rFhd3Z9jx2no6b9Pj4JSwJ2UxxMJKPpG
iSrLI2j1OlF2srSDIo3DvLMDOqbkSbwCTuM9HQ/CTXSirX+Q8P94LdXs3kZw0LS3gQXxculOldXl
/8wKVFRw1nLBSGckO068JykjOVDqMI9SVCB0wO4HoUrwxlF7k8R1gNd/RQnutsxSXPjXhXS6/JWJ
ft0QMpZoKVvXAs6g0X50SAPkG7oXHoUe/wRC1B0DRmvrggI2bbE3e5JiDcuFGp16UREVPoVV3TUU
iwHS7fQ5U4zuX5dIALeCM/lDJHLA6QEPFCeG7yTxp5672S6gh6MGzdh/fCFFsrb7Qu3eRSQRK9Uv
6Y6PM4QGKn2SJYyK9s+Dcv/06wiSdsp6mNq3KQtU3HDGUO1rs6IPcveFcYInGCMYBT2u4VGGNI+l
OgBKYfqkuYMSRxIoqvEkTDq/49whk4fZLZCMBDnmBAI3Iu5i3gjeFqG61qUkKwiH/fxvJLG5205v
dbQJN0KesSfiLUONgUF1cIvNRp55FHswRAq1+eb4VV08/iUi+FDalo0E1utn1++l4s6ZKwT+Ecv6
gP4GZaS6VbHjJJEPVo+YWBb1zd89TQVNjdhv7aThxYiFlrxnRGTGMgUdg7/hpUBXuNS5P95Kt5HO
hL7RbCsxtmsESDtxBmWpre7d2uRjPCwTC8ywYFIvuyJQd1w4ez0Camc8+T+XA/HcsE572XvmAj3K
Di6kAIRqnb/9vSd4IuD+NriKtyqdq2tlgqNcWeaSkk+hUaRSyW036QUL/JAHyESbgoB1HSXK5eiR
/XOM7sl9VTMboF8TC38fTeFk1CnC2pitqonx2lrwxqC5u2oGsMVmyIeuzBrThxAOAC0km3JVE4I9
RJNhvrUzwhKYFHxw4sG7t9xkfbIi31sy8XHNUm9wUfVZXKJs7xx/FkITR+QivtLcwLWYpbtYl6F+
ceU8posfAIQxzZF1405W7dD/GcQuMBc0nw2VaUtiRS4bd+rK3TMXCkQz3WS10jzwpAIZ5vZYdIKf
GIkPVFbTBdy3wtLueti6pK/cxev287BS22hqzMpcUy59VMtaUttruW0NFWvhmoVDDI9QfzFJMILz
++utp7rygX9D9J1n142fmqC0ogIhvxkVoEV9VeoN6+th+bL+S2PaTfJPTGl2oRNOUV4VEfBU+ll8
TE2s0C9XWyzk8YLj/CY9Lsfbqjcsyq7xv0LcQXPU3r5bASLxYbVUG6v31WRySM4rzdm3x+zZmgdO
sOywdECSQGfyzcuV1jLvlZG+KPgLTjhxFfTMJNZifUYYuApuicR5NnKNxhT21W/ZBN2NK8KHw1rM
bTH+jq2rO0Et/aH9iIFpWbDXRRToIGydoWlv92kq1o+ijI+OSTZYKTc4Zk4Xbvt8pmA8p9Z3TMuJ
rPZ+uvpHbuQg2ghJlEBbWcd2PVOJ9gtA2h8G7snPrVMgYEeXnUga/HZrApW3hmRjkkBHojJiostW
FwhPquDCN3+wKojtX5QFNEshxzQOMKKVq+pssysk2YugEh1KY1YBQwWLpRpcQa77ykZlvBriZQXE
/4hHOt5K3oyhWVdAWrPa1yUNQGw00CdnEX27+VmpYlCd+ML8zE3h10qLSKgFd/nV7r/ssA0n9ZTQ
k4jyyZqDqs6xuU3iRz+5APli/XX0f2oCSW2eD/apfN+QkyAes1OdVTBRWnUSAzGkbd2DxYIuvC5n
/XhW0YZMnGhaRuW3JzWF32fGgreGq2ZKpi0KfDtUfTxPzUhg7X0Ihr8D9aL+AF6hKgWD/Nt7jxST
5nbtMn7iWrdj53A8qU5TnIfhM1O9k3KLkpSuYLJaButQgId7hHK3Rr9icuD7SmRtsw1Pz56hfTUm
rmWObI6I5zkr53QNC/u4xp2uCvbxNSB9iEcig5lncexg+DAxubdEoMYOie27kAEBaSpyqNw4L9/J
ySlCBFJY9Fq5fvDHQMi01anLc1jKV/kWFulb5Ey1uUekDEbic+OxoZBOBgqG51+8rWP36+uJ6FV9
QDcwdry0683eTEoxyE4jwQgsxoL00Yi2IChc/YLYg5HgH2riLmzBkRAY+rG4L7ZgD7eaqsWKmvMu
oWmnMcy70Dt0Sp7IzBKUFJLxStLnxCi0STf50Gfu/OBBe4NuA4JT608rTUD8c1zROEzm+zOwtm0H
Pq03ZiFiHEKVNLr9mjpY3hmIfoAscBNANin/g6D+Cdpv7AfLp2bdVVY3Qthxg/PovpYnYnchD28/
red4pFLl8HMfq8izx1GH2yRVMwA5Z16V5AgkQ9+t7zSESv0f4kp2xH1XN1hJFguNVJFN32oKaJux
HaN6jQ2PtvfXy1pkM7kAHC3A734FDTkGUZ7k5Eo3uGvI/Y0rF4K47nqFmPG+M/eZDuIeWH7VVHc9
l1Clwlj1dye3R4Xo416I5ABny7WLR12M02WyGmhhlZ26ry1jpOSxUlYn3Llt3dGrHvrOyHDgnA0m
1hzxL7hZXHHgpcL4s/oRGSVzLWUt14xME5ixn/bktJtVExZ5KpdKDIJwnk3uClXnbkEqg7XQklPe
kvv3GQ/W3VkbE2KYTqXqFjNMXzlihu9HHU4/FNDylqAXJ5Z6XKihczHpVtxWNO2Ri12xMD9J5AcW
h+LlBK9BAAp9qM2KcKiqtrat58nxSv9FTAtcQJTWg0ycqydw6DhOUugeqBwIcAjJ/3a83yKR+5aO
8NlTwHliQdhmf9sUMedvqVDJ9HUKy69V3BkaYpjQlpzf1jcBKiCTtm+vfzXZoyH9ipJXB5/4TpIS
GjjNJCw5SgJ1bw08mK8dCla8XfbBBWlpXqR/HajdtdEK8q9tlbMQERaWaDqTTOgo80m/drNuEvaN
HGVUh7q24DLNSrVXhvDjzdCilGQtSbvJTofFskDRHfp5OKxC8XhCsZXKHgUJujt4iM2cTqr8mKFQ
kjy8pQ/AH6XnL+ZpcOr+Iqb6XjkraugDuWkjFnJ88vkxnK4mI0LGHrLRbPI7HnbaStSnfxY2p5/O
4GYDtxEPobuFcL1vtY1mFLkL859Q3PdZIL9cjRBznmGiIXpyQ5ZLIg5MSofzImaK1BYaQ6MzMmHY
b+ihGmomnrOR928Yri4aUadTAkGcj+XaLsetVlIru1AD8k8L+49xH+Y8HC7ZugQWImBtCbvcSEpJ
I0g0OoclYLLAzhpyvvYlb7E3UrWiXmDUXwkLY6Dx7KplhJ2SYux6vlaXqjHtXW6Zec/khpKbAzw0
Ar+xmd6tRFG6FqoXROtXRrnhEswUnHdnu0md5WLyZRdzfVab49DrE4ACA4QXt+8JZ6Z6qyWNFwVr
wbfRg3ExXmEN2cLygxOweEeBWiQbDDDW2R1TpVIqqbWvykLHQetVlEk1XsC4LW+MUsLwnqm0ZA6k
B1A1pNJOZ8nRyR3pn1bV4mQFMzasq1hnouG0wIFiZdaF1FaOM5+rLnWUPTTlO2MGp0hhsVnWgPkz
mTiWvfKCBRMR8kzrmIXMiGFXOI79guxAra7f+CjPxGyHVjhIB39kkuaE5+gPIztIOvKvcqE1cfef
6L5L2zHKBJ8CgYJcsQxcI+lmAj0O3rR3CmMGOiIRBsMwlkkr9CTYwTgcS/v93tzIq+C/DlcYGXyo
v/bPW9dTRKlVYIpxw2nNkpgCI1Vd486dkaH4q843ymq2IhJthAIfWmvNatsx9RknpGPOiW3t6Mzz
2bCx8sttELIMfDpTvmt0JfW4l1GWssysCalDQbL79BGycxJNYhl+J67lrZvfpDqudwZJg3Bd+OAh
nhwmdQQPlU3HGhAhZkQ2wXB9GnzULdBlB+OVXctyKGxW2RjLQCz8HVklOnSmRe/WgBSPd1vUPr9p
qYjDeBKuhtf3qzvvTcq2OTKg2agB2rnNghq8a2h4uLFIQbNcl2vfw8Z+UwD6L0KJA8Eqfe4uW8XT
VlItDAqVeIcyyPOln1MLOgv0+g9liBNP9v/HuTiOMY6Htxo8XkVScYywdH4G8vh8cLQQY0CWpp4i
7Z3Yl69Cq59N0AwYTWy5GzpKisG5vsGSLO2r8AwjLJzn9MD9uJAC47NhN76mHbt/N9pLQpz9vsqO
iEZiK+M5Lo6Q5CEu+BDbyOCm5c7nYOf4iKj9AoL5hgAoVFx4+TKqGzrJ7cgEzAxVxwS6XhVoMu+p
xm0hJ9XCoFjlswFSmzP65Pz3/HoUnNSLxsYSaP8LpE+DR6vsZlq2DYoMVO+lk7fSZXACjHsPrVvT
cgNLk+bNnqDKHMTGrwI8pvRd/gZjTqm4gqnrlJbiZyEiX+FGRs4GTguku82ahFmZr4jUNxngnV7c
9QAeAtSyo3FjG8m/+DA7152Dd/fpLGM2N6ZJ13ZdvIrGKHFGOnQFnnmQifM3X8a0QSj6k7SQMF4D
fr9PhGi+NEnF0a+Y231WxlnL8oaYwteliGzu5xGSlHGGZR5qPN/OelI0CoN9pKARlU7xsZj1dZZp
EvxiIzlZ2YUgLs8QvoOg/HdyZRtaI+ElDlws5RKX8JQ+5KJdYYNvug7CYFUaABljsbS2bQ2QrjIV
yQN7daNI2muNAaElpWwR59qKdPbJRHLsf31FWT3dQBs0WRtWzzCAImhHpk1MgscAsSblRCrQC80F
wh/rLNusL/SIibjRFsNnavOzGpiuqBxbdZ2tzwUKTo9N7ee/OPDu2HeXTaCTlguR8c7bavPoo68C
IssANxU0suEqMnDpQujRPAnmG/3uqsmbaOu/QJX1WOG3Fg/hpxxYGACCJsD8sHwUxrrV6MphOoIN
VC6R6f5MCpClbfaN2MvV2oZZqDTgkrNBJYfbvUzfL27PfunzFWfuhgET+WgQvl8pc5+8tl4aytGr
jUdMrPSKEUQLw8JEfDuGZCn7+zReRKy82JRVkkX+SjIURAyq4x68+LytfnYONiixyijvhUcEZIog
UmpFoAkw+Y5ec02wTyt7zQAnfoKETDKHglhdCPE4iLq4CMnPagiMjJEMw4r0b/aNNLbKSGGOUFzF
avLJy3fXpqBf0zEGXNfIBMM9aS9jNrZj8dAEVqOdHoRnnWrjyP3r9BUzCMdkqe3ZJTy85R/qxpZj
DrvszT6nd1bHw3tFLzpxOLVk61pIt6rL2oaM712bEIvpQsWcbOryCsbyh70FIbVHFl8zDyaWPnt5
4Giv/2jCbc4YGf6l7z8omn7Caje63kd3xm6YNtYOi/fhQ16V4TcA7bU/rEGT+RPYDMKf1uQCI/WW
3Vb0wFdJ8Ahz+WxZ4+7F3aOvfe5chV6HQ6SAEOKdl1eCzgJZF7Jb96a+2xeAQJJnGRTrdpviM1G/
FDXIGXToodXK6TJKnILE91XCFIscLL1Sq0CMRVKdLF4oqDYdFVWMvEeR5EoNXYG+cn/viDNYG+l9
UJE3GHNQzk1xi8i5SJ+/iZGzoWwrxZqkQ0HvF/wlM/RMuzotZJS4F68gWoctUHcfK1PIVMf1taB+
SGhUJHNYXCXnsU/XWYNj49oLE8XHEgCbqMTee5ZhNUm9AzOYuG+dIQyBItb7Niee/9VDCvoTncXH
g3llrzJLKgBwjkHYW7h8kHaEFa5mrvV23p0+X7SuzTmkqu3UQfwElLVnGxFz46XSzGpFePQP4ffo
vww09+FywvLlcp0nGIF7x1WJ8xYxcN3ksAhaFwN8NVX+EavVrG+UDUERyWYnbfbHf2naKJLp+MQw
M9C2pOdLil2YSnLql6VZCo5cbWZ+hLX2mwqBZ9w0SGLZTYWuzR4lMNA4l8AOW9D1178uJS3Af+4O
ZarlzChhUe0xfJXm092BIHRVbU/p3JYcSBfKUX/hLXLY9G8PTpTjFbEDw/jUU/ODC5IpcAZaGuPL
gbs2ZRkX85550uVRQUDx92mX3X+Ck4jGWZtYdPPe5RJVc2qwaiLYcywZDlWFUNOSo2Zdl6Qgsr42
sZ2pJ26FMeJw0LbiON4Z2thtXFGZBdBhJOQwBmzyp92nwp3Bc45Q6HLCWUU3UBhfjysp+Q0ISGeg
rWYpkyGmsh8Qy2ckFXPyBmd8dkLWEeqhGvBITSiCPIlwAhTaWC83tJ0EGAOH3l0IQy1IuvInOfTr
No4GLH/4xNXWM8b8WFhvzgL9ippsRQrSnGg4qE4ImXBq2bUj+DKDMnL21nksNmSReyS4Exx/ycvg
kOSUSkvVbMa38nYogaZ4MQrLs80dJQZCSyMHlB8MYXJy2AT5c6hsWKZedN2sY/gGQwB2/2Meh6Po
tpasjuB1lrt47Bw+lT2M6vfYurJRhVioTsdJQXxK3aG7GYwLY1V2akTjdcnlbsC0wW6kMfzOKWM1
AjGyYQqiLH9MRzyQ/w6KvUki/lk2SApegWd38si1Eos7JUCo/cGuNGE9NjNJ2B3sQpmOXhe/OKCx
Rq1ydM+XWIlJThpsVmyC2iyKkT1puL3aExEwdeh3bwkfz5nYYHTGpCZZMfvQjJc1LoK0MGaWK+IL
f7xyR+DkLk8ZsqJ+QeB+F5mS30hjagVJabNLa47ga4jJnZwNUGlWQrZO4hoSfrBmcKYjgQ4npRC3
Cdr0W6706DZZhBIys9GpeDakOnBF5LIpGFib4Q8gtP4qw0Xe+acZD2XMD0ew1kQDzCNdjJCe5s+0
g8dmKVbDrhvPVYbPekXH1Acntf5flIp11YgKKGPMj/2plDSC1OT6ea2fIi91XrQc4PYVl5vKf5+Z
cXv2e9TTlxEIpwEDNxy19zBYp9wuCcnNsGbh/swN2uCCKUWmynCf0UQQC7zB9jTavhEVBoobdj43
l9BV3gWImC5L4Pzh8jBstDn/r6jKcLef5iBbRrO6NcOrBlNAnEPkEMBE6ZtJmRSca5Zw8EQU8l7e
Mdf04LIUzxnGyvJyYtd2/vbwKIGJ65ToXoTJTA9WaPGOPMTMjjOcsTSvCaWQ448aY/Ko2s/tQTHF
wvJGuP8ZIgNi6XbkixTfswOcQJR3BAhV6Nd7dnCTnWC6ETvtkbub6mTUznwOcpZ30V9BGH7pj3p3
59YHNgihsFzdEqLLlsKO5wpjCHTITTClPu4kU+nklFLW+oSfEKMRdhk4KgrHPzyVzGmZ6VHllsuy
9FHJfObdv02uZ40tbYO1MelMBPcio9KXSNWPSydbivQLOMLoy01yJmoBwlmEYfA2FWt5yECXfl38
etDCUr8xVI5BlPaSVa8G3h31B+rGNFDufzEww3gL/jLFW/q3uu47uMHoQ55nHWN4yvWgKMCHEr3A
G3p9x92TX73Dc+rC38Mm+kDaqvJKkUuZcx7eSvseO9033eQjCp6u+yRd0RYoGabQFWibRsvhwosB
vc7mJMe7Uer4gN/YrSLhONBIyWvSIfebZCNFw1XupdbZp8WxAZ5pjKDcJe9kDAcZeDxc9J/PecIZ
dUoSekFhXSLZD68m4F31g0xBfe+1zcilFwRnETzGNkfKlAgOvZ11bhSQFYfSJyQWC8b7vCfMn6wl
Dd5q8MKvgX/92DxnTMm7VRK9Puf7hbjixzL0VAJM6N2Kan6OlS6flo+3N6TW3KNUJCe8vJB/7lnx
f3gv8J8i6lFHl/MIANXYwJ9HRxncChYS1j01Y+aFBDBd7G93hQrEO70pETXHpfvzffvUUgXpQwv5
7PQbA8SpxnvCF43tWMwrktpCsCM9o4xuFdCKwa8y1O+iTIxVmrxTH9I6DKSAfGn20cOGCxYLt6y2
7acJo+ueS8tZ05DMi3dcbrNXbdsAAI7wGlusA1OEyJerE41jneCNaqXOS5/9E6rR8dwJZE+2XrOd
z8qWrgMeELbFxGMNIE5gPMujJv5g8+VibunwA1E9whD1ex8CLV9vn4x2uG2hCX22ht8/8lZVyMzi
lNvfV59JO/E5kZEPJbIAoS5zNL9CIEblqgH4yqhO3Wneg7Ek0T4p7Cd2lCZTGS0UdBfibJQu9zkW
SMFQTldXru/zbMnDvWwZ9bK1LwCXInEubtfNdyFJNNV/JqmZpKOSe6623mZ/q31LS+Fzi1+CLrnm
HUaa70LxvTo1S0E4BWXdhKgk4NDn9AN0Ya4KfqeRK4hlpwYk6LS8Y4c0UPvAQBoXOgmlEInZOtNP
G/4HdxhUGRU/igCtFBEiPWPh4FPPaAGWr9cvxm/F8ECLlGMl46IzLJs1gnfuaiOrujLY7byIejfO
u36totq4LWmwBfOuTE9lgSQKYnT5IuyDOy/u4D/tW7wiA5vtlVf7R0Fay33aLSv1U/4+scTNQOe9
AMs4gsVLHHu39YItXjPNqxbPsiSXsAWFlAqiIfGr7mqHRvWid0xc/o8+0prsJEYuV6wpWxyNgD8l
PQDcBUZc27zr8U8dBWfMdyqPOkXCIewqhpHRIngZJXDx3F6aYzv9wel4ymlWW2/rQERJBwEpRSsv
wniLIGRqbS0tQ1BeakRA0lJZ4Toum49KXUKQGlos2/Irri3CcyVVMFWS3+wMU8Sxl8TY2paZcRyo
FeeUPAJ4wa94UYKwyN5WzakpNZua65qup7TthdjO2p8xdVKAijCq2/0LrpBPgodfVX4+AizHSJ/j
WxHKo0vpE3uH2SIMTj/DvR/rvHsxVe88qAtvoS3r3FmtjTvcbQWPLmwy6lPGDySLZ4VBaxqn27sZ
WVk+auFndAd8mYOQJixakc+JpI/sSi8ZULSC6XEEXWp2IpovCNi7noZ8XrwfRr/kPqRn6JiGAuJQ
VJnj4L0zbJwMQe1mJmeIZsgJOC36uXPOFwBQ/h5bZltvolaoGXEteur4koBYm54WYL5wl8F2Raed
+zwGtAj4vEFemRhqlsDFOoHGGxEjCbpMXcBwqSHIovWlnmujGq8Q/bdcecDmAl6Xx7cxbTmYRWAE
bBLTlZ4h1Y34mbj0/HL3BkC1n3ZS8awIXhhetIRfZBWbKddFsgyfEYzjvHazY+HrjwBxfvEDcpRY
cB4Jzpj4Hx6akyKn3TUMuTHeOQlC7o6krRe063sJwlF0h96jEMUtMjGx7a7MQTFU+ptPT1SyJ+TA
OFbkBZdlKzTRLoh/JOTQyvApwAyOZ0ilCN+al+ZGGJ0Ljb5riG9wDEedHPgiw3BtjmrHWnXg0XDD
5rljVpPdJ3ugiYYkN6JRRvcfIZXYD6N1MSS92GAfdyiX+/2W7NbSxcV6dwRsd8vpWnlK7Wfn5Z6h
fYdNF5hBLsCFMmTUCtt+dsALY/XnAejrUyKJiWbdOHiIWOly85H+CYqM9/0ccsSoCjrSrYk9RFxy
mNVEUiAoIrl64AQy9fIqu9MfbhTb4AAJ1W6qXFntlFYh+JwIn5Pll7LDnyc6gE7G40ogsb72yjNa
2K2pRdsFXOTtC/U0qwGft3VBH5bCk9xgRASeWtyryxOMjeplr6QKKeSx/iI2LzOPppKnO6MjkKPe
WOrlsaEW4czWmftUfhietiWV5GZ6YDQzowrtiQqAc1OFYYphG3V6g8lKVvmwV6BcHjKRye6JcU55
fwCHilI8LlfZtx9px3tbGNYtKttQ4+liBt0szX+13bsjS16qqhAmodu9SZJGB8Tq4k4EhhITW86X
MuGW1bYEjAKFMGjZbCpUa3UvWQ2ZfBOvPFWhtLHDTPno+0oUvoqsITCia6cnJB1f/BhSZap/dTVA
nzv0ZH1khzs35oOuGOT/NTy6yTwZOSOyzYPTF0g9Wrd3SUs2TCAMr5uf6Jj5FK+bT4RV+ZyAD3yV
dzZQJ0VFdErzDdUQwBLCru61mRrmkDZYQz+9PHdlvAe01ftQqKEiJ+6fLE8xMmfmbAtanDk/c6tg
YVVXfdVnn4HtEsuPRi3GJmg7si24ujJoi5KuLkw1tMa7czB/zGdylXL9oMgmbX73N9O8HI5nqHzU
ElB7+u0hFMYgp32LHyTbJowM19fLjY8m0UdwnAAaGoprvDEnWxJoji/M1ZCLwOuvivruCOTnr9PM
+SjBSAWv3wJoCtXi1LngV61/WUiY2D1StYqFOhFtWOXF+SEcefW9BbxB45EO1wfcmbr5OyJP2iDS
VPmCD+SZym7Vb1qmuASEJytZEp3mdrGQigfJO7glIXsom+78PEn5yE3K612vh4YGZl5fAHs74nNM
4yrrr1tiioUiY6kZ5/OWqsf/jUdxWdu3UK4sv5hSlieijXPbLLiBbGOzYoeV3pU+pUL4hZPwihyd
lIkWTw78+t2ZqZokRtsLhnaA+oLMho7HhG+9Mkv8PrRYst1Qi8D+MSNtXNNzJkyDiHV7ZD8ISs/O
qaeN8rc89GmLGJfDdqESpND8Cvp+y+smUZ8kkHDkLbOC86DFvSRP1qyFctQIyHD/keDAN3iRdgTM
tkVhzYijEAdaBwtsrBBA1NGe3k3Ad60Cc7fZrFomiiHVmyrM1BsxsRVrq7t0wvFWsLts7bl/EW+j
1Fo2SCHEIigkzi2ijvKWJ80qMedM2d4jCwiWqJf1JP44W0/i64sb3XtfsmDdr/aUkaFO+AEa24xX
Avdo+V/8c6Qvbmq3Z5WngUBDorE9UxIbmxArKKo0NE54+6BdnybZWOSHUzKfe3ryMAFC0KH15fx/
KW45+TZpJKV8NLLaXJ8VZUQIGDgorLPrpj8XX/Fs17LRDmfEUn6frB8Y87E+dWn9WxqEKFj+VLaJ
Nkgd6URZ4WXJm88YzJA/B5wd+He/kqp6z5DS8MXkGqtC39FaWcXF8xA9t8WpktG64Kjw6qWKJVTO
/PGjNd7Ju/tBhOWlw0eOcjlUGo+n6D770inaD/0u+KbsefKTOJuxY3eF56GDwsySrdrrJi2rFSQQ
VOt6a69jPH5xlIJmPG7wiimC7XLhnBBzb3q9WZXCm+zfEABTx92c2XiOCPrVdWjqstSQTeeldqsi
2o3notlMlBBWZXoAG2Lcu/9t5HzTSLxJ9xPr9xj4kXrEHXPNbaOXFk9NYSfifLwAUdk2Su3z6Oau
njZ+W259yMJVa7S2R1cOmBsZJleGPzYS8g6R7DFjTjaRRe1nJlDKMyfYmJqLl93sxtpQ9OXqbR8T
T2vt7H6Entizr+nh2/wsKzD03YGIW9JXw88V+P2bRh3A6rMbdCR7uNVHpQg1zkspqLamjKcXveLu
kaiizah2J3ez/DRKisQGimMyY7vAjqyHUTXeMSD4LR0dQliNoPH8pvPzo4IUWor5tVQr05RM2T3d
ajRyS5CSnlEJcbCu2op7ItEoxtO4D85OPpiIynnl3jWRONBjpUGIfCbhUNRB0bUEog8LU4uFKvaW
fu+HIRPfihGvaxyDYtViA8Ovdu2GNkVnk7vQaQwMrUjxOj6HuisVZ78wV8FI35EWOeEe7uNNz8+k
HGGBNVavbnGbMrV+l8iEM33OcaZrtZ3up9D0UxRoqvO/hj1F2l76IYjiFe+GYLA6XJas4i5SQ73H
SwNmC+Wg0DfV32C7jvtgAp+qVarzAeKRXI5FYLm6gAtKH2h7tt4BnEcnMho23R6Rnpbeb8dQ8J4g
xm7lG7dDSqjLlfW3uijmbC5beRROf9bOOGICb8wRDwQURr1X0eAio+h+3eRQsIf20FurJTKVlltK
QzPdrCR6mRbkLzevNxv20258EtnEl4UbBoBI1DlmRglH9oMguP/gIAdoyziP+Jrt0GuHdoJFeUMu
Lo5PUboJ3Ns+1XMmkNNFuNzl4coZ79a9xg9xrTX4fXYmJ69EDamFP81w8xcPc2/F9uEB32O2lb/s
hlOg6Y4Lnrh3NPUJKgZOsDBuXY9u+BJPofqgSfYP265PbabRQ7u12l/yRjzb2bSe+CCMYQjZVGSB
z1EyIT6TAUqYLhTptvGHldBaL63OOZQfTv/b5kNE1J2L6NeWyXtMnpapaSUANehIULeTGv0XduHr
Uup8699eMBUJLsBQCFpHfaRNGlDAIWI9bYdENftjgNxDL/yTAfzcmJA2v6FgsDteboFx2L56/36S
p9ZlX9SxzGRgvx8rxzsiWMObp+FiZsOA2S0gBjUHWXW8HJduEypHjXXgFf3Ho8l6GC31vzMe+AW7
xYgOq+48yQA4kqmszzpe0M/rMWbc04UMBpwm6QUwVRoENalUZyauMl9A1HQJ+vHA5XjTl2AHZ/j9
6RmwQc/x3JUBOcJJ5K9+iZd51bIgLY4lHYJOmOV7sVc6Xa9V7pe9zHykMhuLAlAFifuiNvs4BTcW
kuqxfk5s73aeU+5ARlH5OOiIFWJ8ojNrDa1hNvDhgo9Ln0r4jmmBS6QCCVDtVkBT1tgkUQPEKdg+
Ee42gphL+QF6DfHGfqF/RaJf5GWxX8E9vHAiH0qcKZXeYWM7B6JH5l9mMILDH19bEVkRoc+XR4fZ
dOHLJ5OloJ/J5+vJ1KX/JLMPqmLWEfN7VbVh2mlwZHaJC0evzft8gu4Ap8EnuvHmG9IrothtOeDp
BAY9zRR0dPIk11Arl0lWVAKE+dydPkO5SluGhPGAYDsLV//hLSW6YZLDLIMwZi0xpsb/lduqxDxB
1Sv0n+dhh74a0h8+v2VnwTu7UbNOoQOGW57GBJ3HO4xrSuiv8hRVa8rbpRNEeaQey+eUXqi2ZxVV
5xGR3dzDZR/PbNE88ADhuwNRpRt2tewqgr1UJiSjOaOJe/oKiarm/WUIcZFpi6oB9ybaK0N3Udhg
zq8KELBgVSDKIHsXOcTWcp757X0i5lzVlddT+cyL5C0Sm6SeafejbjCyK4osxtNfZadW8TXNskWp
3TXW1MGnC42PBuQx3o6yENU3gy4u6MIPs/1IOU/ceaOElrNy6mGfQxxrZ7s1/cTm6lW7L66jGrE0
PO2z9WHBvZU/pwKL8rC4589o0liYGBTV5UP1qhsuU6C+zcJCFZmUh09Vq5HN1PspKYyuNSAJot0D
dOXMZbNtK+M76joN20Ciz5gTbwZqFyyQd60G4SADPoxPvWLDnpCfqfkhyf8LITS0ydBCwmnr3mlP
Z8vVRaSfp73I75BhPU7Hg3mI3natC0+IcWnjxea072iVvVhOsFHXA1aqpvkQRHWy2yzaKwA53yQD
emaGLegY0fd2vU/VWwLowV9ZIJXxEuZkn5UahkCjta27igfElajKlQ3/wB0/F73e7ioMkWNFOytF
hxZAiBg+4AN1IO6Q4jrXN4PLhsJIjJpaG6PY8Wrfwt8KR9Xtomna2AG3UOvkfkRSw7ZitSH1GgrF
qomlCUbjeC4aBVXgVcaosF/RM1o1fPSmNFe4YyNAxxhEi7E494eUdUmDX3a/y/0H3qRFNn+1gYPA
nInBVz6ufvZuywyKx3SnGtJAJk+6mBJZKSvEUhxZfDqaRxBmTjHZdbHUNttkGX/9gfKEFnYrN4rc
LxBUUQZqqcULRZE82gQT/YXCSb1hUGRdwyov7izXhjPniYaYwSdpL/B4e8aN7Ehc+O7R1ZPsmWpJ
9V9rWP7QIZuYqnBWMrdZfGHv0nPHfQ5CuEDhV3yJ4RM66stWLIQIENo4tfesqQbYLHz4JwUjoYOf
gnQsGQQFZhd8XsluejSuH2c3oBXxCIYbQ1PZIUKqWVAr2MV44WrERjp1OhFQz9HrDNUdYMpCkvKV
ryyKzUspTWzzhBWtzBk3qp14wzyOL3QaLaIWOXBy8Mlce0V+KSRAJvGbWOsPOfpGvf50YlJcVuPL
EWooPspe2JgLc8xD8LoBpraasI1DhfAXjSOTxhMwlECFuLWY47kU/N+hM57lfS02xxE5ctmKhEjP
wiCUCZtkbQOe2uztmPPFmTvJI95J87Gj5Ll9OZSq7gS6YFmfbE3ZW4yKYb5NnTSfFo2xJzGtvn7C
UVHhuyJJSqyGg9EI4uTfrVIIM5q42IAKab5pzo0YLqFrwmGdwwOxuKgfaeWA+dWA5SM+hiSi0BUu
M4rb3sYQNfxZKJVddfBXX3nHpLt9AFzpqbxpaPcmtyzOUfMYsYyHI/lUq2NSzG7QpIsK9HOsOzGc
yLwETUsnl386oKmpEhzl9RsS6UymjN1TlaGZ2N+fJGk4uN+g2h2jxYaEv6XCTdd8f19v5BuzGl60
0D6QyEXcJZdztyTvUER2NDayxkAW+Bg19wLpTltsHGcbpCwIXxCzKEICIFKhqIr5ERWhORa7VvlV
NfSiUeRn688BxPiKycqG01Zjh5DsZs4TGxEG/hbBRXSrYhckBDx/NJTJ6tTSCu6NTWrW5giEp97C
9LATeR/ZGTTfJgB4rnG/r/Fq9qlDJFKseFc7hQdh1IT3ZvsirdtWB8qrDt3cNc7mwnp3WPCOq0Rt
zxmm1/2hJVDkx7OFC+6y2nhYA0ujp8r0ilW2U/G4fc7+pzfW67ksMrJK/x9sSydCi2hUxXWM13/I
FrDRh1x6bxXC3ZnqDKPp1YU8yKYu5z3XxPnEfUAZMYiqd0Yhy8WA5PtgfCBSA38QPmU9bg6IUE3N
dhaV432di7Cv/d2AI7Ue/1RT3BcH7GG9OwHE63CkOVXxNwR3vVDs6QW3r7QvvHxnT18KRV3rRdpN
70v0kR5bB0wC+wskVt9inWcy8CxUlRPK/q4OalR/i1PfgMQ8B/BX+A6mHpdEasKPWJF8udyqWEL0
YtPgLkLUNvfE5yqmzFSC5uMgA65UhZgm2BA2dQXa8vEiu2qvSSumEszEa97CtFmc7GhbkHnMGo12
VuHMmnY6tNxl7YsSGVWXWG+jTF18Ous9tfE/GFymu3iA+gdsOEZddOBOPqPsJPPRalRSqthhUXBB
OkY//l4bWPgL6RPh3HxxQvOEWDTdepJsKzTDxNe7YeCRzidPfW6f3azrc4nAmPZx4uZTPMTs/H59
LmxJArmjlXRb5ChPPpG8jQ56g44BRWAZpj5rDqPQDx6tphyG9YR6shds5ES3hsjxgv1ufE5gEGfN
9R5Ge1fW+Q8bcyo3XCPqm7pg+oFOrE5kqNAfS0TQm5MLB42yvLGi+9ocyRZZX2Gii26yruRNPNeh
vph4QHyUsl0JZBpIztw/4xOfFHH0CGtQIeBf3dF6VIqLlHdsCzZXlHeE5taLVgQJK4wNPD25/oVu
GZ74OEa4Cxn82UABaf3fEfujXz3LWxT45rPTHKXf6pU8lUTwS+j8NQ4bp+BFaa1aqgon9zPGA5Oh
eTsqRUuBoPONiwjFMZt8F3c3NkF8KqALnO3ActG/4pBqM6IrLJ2HOhvz9C+Xs0YFGqcIJ14DSjXm
NqI5pnK9VVnbDLE22Xdl0305YyLeaA6gxG6/gAkOa4H9Bex8fm1Bw/owpWvprnyAXWB5Ok3Y0tAG
vilUIgge+FvgrnecAo7pwvvtJJVsy2DBc7qUzn2rPeo3eyRLSSv1XmOgcWTM6rNRVxooPUWlUvQV
fEdA0o0d7vgEK7eWd0F+c2iaAiwK8kviEUGSVJbjx7db+QDeRNWTBZ5kCWlv6nGI2teFmYEtzvLK
Sc9E/pzsNWPGz6bU1j3ooVq+b5Am+brEhRRnh9FdiAR+Ix2KN5/Ed+gNROL3ePI6FLe06tFOK9vY
+g+sEX3hhsAy+O1dfWIcuIGipoe6pqq9klnHnwCjj35Vev/zxpIGTG7nu6I30uoIwzaGt9w15ch8
fWx511G0qFeCa5shaTsgPhA0UEhjIBpcWPO065THzHDi30RKltOvRXBiGVSYmw9d6F30F8z4lfN+
pGDWZyH6/WPlwPmKP86IR0f6fNm+jJE3wcSpy53b11eeAbXfrHeUBVgWq2yDo/jK0i1WtfMpXBek
/IeD8aTqmrOWi01y0bA2qvoFJhd2ZipgLOw+VyPOahvApT2LMCp+BHr8hl0GoYmPvmZEG01M9n9f
DpmUopFOgVEgc+MRHl3YFV2nP+XxaMx8emtXEbzywjzKbPc6K3UODlveq4vJPsQUOk05ZjDZpadQ
sME/lCq9YyF/8LF2nARylqyYfQCe9dhYy8y9rlQZaHkcC/rDZ+F7BIS640Cxc4KlX4XdBoj3d7g9
77usdhUtuiDbNAEL5hJUWT1lisyQlduKELQZS835GYKLw/mYMZcM7U5lMM5/rQXobZuW4AvIhBW5
ZZSNpW2P0BIC4saqpENnLvZbiTZxPSQFlIbmG905IYT3YLId33i4riulSd5QDQ6c4PCGM9XOeXAA
15pvhWcIP5rL2FS/Ad+6GlLaUYQdy5C4a1SUIsInIujiLJGp7ec8b5GIsaHtQyME8UhXWoPvkNin
4jOV7YUXQRn5IxkiNeFwdwOf4UjXi/ovz3RzUcKBGOUn+frF+CJGKMZDXaFVZnY94T3zTwRcjhtc
oK6hPt8hxYWFfY0AxWoPgSoygRfAu0UPWLYywzFh/pYAnQvohrkwIl3jAit5WTiETivD3jZ0rAni
/fzpHflS4M4jJetjWOw1ITME5vabja37c/bzDuCtsp0XYD+ZhTSpxJd7pSZN6R+viYJFSqyy3nX/
RHQGS6uT8xzZsj+4VtsRpjE3XixGckhAbKglfEptELcA2pHrc0icz3zgGNftxc/sxoMQ7y3CGTFy
QgKA3UxMYLN3uOREjxkvbyvaigjpTNPk8jupHkQ6kfqXGCxsojoKgHycE5RsSThFQlJEvW9tZoAb
6v3A/8ufFIL0WbA7HF3Ced3OS2g1eRiGM1J/1ubsooRnL3nrSuq+Z+yiVGZow04Qhjqe9RbA3ajC
LUHpCyViwI1whUL8l5FwyZL3ow6BI8qeEaxAbZ50Jz0CqcGYkKHGgBoBBhmwLl628XsVLvBd9eQl
erghUgvS90OxcGJ5l5dMsiEjm+3DV2ltiFXldCSxcU6B0TRBlxe7XyfZb+Vtj1yZ9zFTzlqj69R8
eiVrN1UOd6iRHxdEN7VhiGcpiMPYnXrKzgqv1Po2Q1THk+dDhiqDiFdOAw/Vdt7iidvQ8neMe9Mh
No3qs4eRysFdDFWeLHKHJ3zzLHiQfXNw+tXgJee4w3k0ptE8UEoOPsBGy2ecKuTDOfoto3vYqem+
mjzXUrXfG3i7SBr3K2uZL6gc7FpNLqguDfEdtgsMVlmNfwbSKsk/uNobTQN7YquUZ9XILZ3DGi5K
VrihAK/Ce7XuGARImDAVAt3gGoyATF6VM4+Eg4GFaCLHMMiB/poK+ZozvV5iEixTrZ7jqP4VA37H
S6ewaFu7eQhN7zdMfpXGU6JbnT80moK+Gj+AynA2wiwooSETyl4vzA5h4krnWMwZTkcfpSGxngIU
l7jw1YAmBhM2dXF5VO6TPjj9PfmmKZIq0D2SOyRbpiFP38bpM761hv40oY/2gxk1PobnPNzcnXWa
wGsBhDaFhE7g5MY8+qxVJH84PZZMj9EigSCAQjO6ham0h9s6PECKACaBZG5tGnSs4u61z8h2Ro91
/T0qoRLiGxNb9Y+9MBtpDrc8/Amx7VnxPS/yP/VQ1v2EhMIUgtSdo2gXaBY4HorSc0GphZ/mbg8m
M4jBCcXzgmYP2pYD6vR8zjADiLm4WOQlOnn+OtyHW3sOMMypA3d4qKGuSaahxvdNXUgtN1Ww0zI1
v2iGwwAkVFhY1lY/EAgBgL+k3VQLo9CDtv3RLx01ccaUfTyhG6dq5c7ierNCjABCAwP3ScrMqQd4
eqwAhTPEfl/JT8Gvc7IXnBPYTITvuPwkgy1upWxzjIg9pcNEANaMvcna3lOPjgOfmRlSVoQo03iP
EQ+2x1ppH6mLGnPYX9BA3s4kv1Cz3+oRgMZ81KTMSgyOgBPBhnoeVHUduDQOp6FmVVV4TwobQS2h
mC61mgpIJtj77FAlixJK+3KBQe6LxSf86Nd8/CSVkJNtLaSLN86SotkjzqIC89LXE47jI+nSNwam
KAruperMYMud+6OiWE6QTklaWD4YXjT+oIIyABzH9Idx3/6a3+y1HbxUnP5d5IAKzrY++5M45cLi
AKZeID6CRMdVvE8u22nWGK2C9CdCN60bkmU/JFBWbvIzCIS3yu7A9HUOT+L8yKZ+LT2mauHC/mPN
nW3Dd1t3EJVmvpKtKAUSSWWGxawkqp1xmkRC3rEUXFgIs3X2RpDEbNxYFP0MA6FarYFDMPHI7oHA
E6H1adrHEK35fVYGHmMdQoZapWucRA73DmYAPdOvUHEUFYiGMGc0fAKr/CBlXwfuL0qAkCr39tAs
2sp9mq2N89kPTY7M76HZxWMwcKz7jp2LL7B76TfUthg0MVYHWTIhtB4bm0xf/q8RncJmD2bnrCOW
OKclnkSsD3eHqozpeASfELctI+tTtb0K6rJIZbuz+Yk7hVkWJpDsIDuOi7zgTpBPQ4HRX7vbCa/a
OAigU/jOH25dZuHfcBKEjpMjnntUBmjmv88fX8SjtZD1jrHoJs16FGMH1kif4SzouSo68xn92FkO
AngAGuKcyeOxivJnmyr+94g1OvpfCtHLn7jxEdQPuLqBJ3aRjdyBksj1O5JV1OVGmL6Z8nsy8vTE
F4SRNkyI5y+qHZw+eTxFgg8F2ORdq1dDIc2hVVh2lsYPMYiRdkM+oLVLFWbV4MdsoBld24HvQ0p5
9cOJxMlyvGm6gIg9MxGBjCMosZ4w6Jz/wGbeKfgIq1KU2kEJRee0gD7QBZ+75UpIOHYxUtQIJsz7
xl5Ot9XQx72MrCG50uXA5WqoebDzUmIJJPiAFHy8DEf6XOyB0s1t100+fKfqj8F2nj2e7+GXAhBl
HixPeAeR1VccSUYOdXpX392i6NVb6Xz9eQq3spOUQD0rybyAhQxBeWjKw4DlByzD/JU3mcu7+zBG
OjC9xetE8pghfsVB88oKcgLLdedckzXSLtENKxqIv2DApyR9EZp3d0aaQDDFpAkKV+QVFWN7HwgX
s0Ht4LhU/iRT4521Dd9ECIxYTqLtadN9Lj3/OJwU8nEryyC8jfwZy/VI6PgpS3op6OZBid3Io8D4
01lMzikuK6mEwhbIPK9fakHQrXNANGcwyX2j5Ncu4XsxOQRRPJIOqb/4Jr07UylmsVUSwLPPUFb/
xTAPM2K+W4wRGljtIHUR59mbAarrmQKTTkv3SbzQSyyoVVkQiyt5/H2hM9qne0rlZB08ZxhK/hl9
F8KcP/e2SFkBnHk+/6E1/XPt6TdjkOQb4NNXV8BpnmeU6QvPzQyI8Pa4txMZEUWaq6Ncm0kaPQh6
x9G0uNr0D2Wg1EjSYuQGRPyrCqL4Pl+yrHFjUnmvV/GFFz149vmu0W/HcRjj6aFyE5wSHt6jrbMV
7DOJUl32YVQG0WFwWcGFHSTP7y21Gkco5U0hD4LPOfHwGjb3JlkBduBYgJ+8moWW69Up4zdO3JtW
5jy0pBi3iDKAQIQ6/W/mXuipnCsMWMRD8G2BU+ctI731re6eFkT3BTEKCHKTb/dXoo07dr/OkJi2
lu/Nh7DkXyFjQvLUqyUDCRzfGtzMegHUbjK06nmLZwmJH3sFfIIt+++RYbckOp4p45i46MY8s6yr
LynglvcQtRUmJw9ebtKAGbrowslYZkdUG3s8jbntm3oCrmAAVZoT+urDVpRHDvSYBMBE0YEvT2Cj
qU2EznbyG+grybqAOnMJYpWm9HycqEG/CgQuEZB1I0BNTle+6r5p1AYdjo8LriPwo+KgBnNVYapz
aDr9BjsBuK4GmR0NscQ+T4LpUAcNdunFurjlYTxJwy1N5pxBacvIhHxC/wJqeVh1VbVTMP3NwjBD
CuJp49GbYiHqYyrmguDVFrpHjuldgTWN6r9E674jC0obxZpRfk+zKePVpdlPJgLfVVVILB/xnEA3
bpgG4yFzD7bRfakTB0TWznv96hT7kJscPxRo7RnLSNYInb5zSg3acqd1HJvCaWSFWE8Jsu0eZcvm
p+ASErUfuRwMtnD+A11A9K8STMdSktei1BmqNPA4hDyjZNPSEoDRw6UqaRxuhcufzbGFi2Eisxg8
HjbkULx7EuVIbBYB3L6sl4EkIedSVtsqRfcmNHKpmXlU4XWYwMUGQrvztPp5t+03B+tJuoqXY3BI
+Xa1zmcuiPGj/6Rq76rmnaidrdnKG325pabWy+b1Z6YLQxn4Q6Q3OTa38QfdnNcAYcO/09tBcTWn
eSY6eTDCraek1ab4fW0VqOjnpnwVBd+Svu0oVFsp/8XNXtuarSyZFCExSUQVVktyLCrTAZnmZRbm
WKWBadwCchX0ARnONcfYYz9xrObCFPzCfw5uqo9ddpI7juyfbez2B7TJhamxhp9oS/GB4tp/+s3J
IILDX+96SUxFvm/OhrlEsJNoV84QCllj7DdZcaaTjowsBIA6XSVeAIT7SplXlB1Hb+iSrvYgJ2Yl
sac5raOjaFDqF9U1S4hDQFu12s4gO7Ly8ePFXb9lhcEmfERz/4uzCyEIk30Y7Dx3iYZOfNlPu+7M
fsMAEUBqebKE+qmWgI+Fgh6m+qJaeRfLfKAzbXgmKaY5uced/Wdsoiot7xuNrlPB0E/RiUW/UMP+
UHtDMy8ayb6jUxpDUslNDHGUzKGU2ql3AsawnAQWumygMFzbtKRkxo0HPksZG14BviLvJSiOQ/1Y
SuabLIkz2OOcghgowtbjWZQWVnJC4xv6KBsFYDKp3bqdEMJxv35a4Vw3YpsM50mdtIGpLiHRxt7c
iIXP5Pb9CnkXhQc9/xhK6JH6K1L0eqV899uWWFu0p2xuFweOuqdWHoeI8Lh7oromqVWV3XF0XiPu
0OdaXSixDhCW3TqLxv0HFSUB9ENbgvsJPmQBsl6+Sv/Dio9fhNBfGEgkHGuoBRgxDbzwCEveMjoa
UK/+0hMM7gZCXPVxaCnVGM3er9VZdGHhOsYPRi0XrIc7oLPFK81nmf5VDYtTExQVXk/UVREtXCPY
WtNQ5AOUfgghXhPJdvUQ/MBZF8LQo08ZrhwjSs4Jd5s6RPmvVvs/yTETEHzpSZP/IpBwFSaVEiaF
KAXFYth1Ktxu/oUMeaxkBuh8MGej5B83jTFZ2H0GqHw5ydgHTLMUK4hlM3WPv43m9HDDexZSZ3fL
aC7+4nk/uJl+j5Yr9LVGSQYAlhBqzZJ8UMskeQU2Gj72ABT0MhIHGfb6dOdrfc0JFmn1e3vTc7Ev
UZ1KFARJ7tR64Y4DR0r47xwXMReWiYC2uC/MfHCtyJO2cW774Khs/Bz8v0VHgKr66NTNA2+BoudG
xJHrdFyncUFpsJ+6j+3I0O3rVFzaVqJRuEdfszCLkCpF0FWRwAe4pQWBEJxGLaIWLPyfm90gx+cE
oJhYPy5TL9vWkuZzKAMKJnkURCsQ8/AZD0slm+Zo5PwzoiJ6i4b+cGK1ZNKNS9nommzSLYCR1w5x
DCoIn4S/IpVSre4x7FM9TIt464yievevoJ17b4lJao0tpf/V3AI38TnFeCA0GPi+311ngz3+ApEQ
RzFs7X8Z7VGIyz0iPqY+KP+CbBpKtob4zLQGs8p5Dun9dudvjHSXKul/W6vmwQjL/8aIsT2KX5nq
lvVkV+yUGcU6AreptKq2yo0D/Fr151XD3rD2kAnUNwUrozP9XmjAzqxiq6C1B3yqAIQmqJFaOP2i
eMdT/lNubQX7vU+NEL1ljwa1ev4tdIXUZdcxIDeflGiDFaW/QsW1ZA5r70sMW3txY7Nn7derKMqz
ivBUu+rHXukY7ryHlNPZjbwXL9E3G5aMfmr4pt8T1FxGDFr3Q3vEzhmw2xDUXkMB9f+hiVdQR4Lb
s8kVpb4Hhq5YlnC+5ZNupR95nuNJzQb1vaqpUK/jRt0BjAP1xz7aa94mApBPkGrCKHKQVzcakrNT
qGQEg0wdTLzdgww3Ojbm5p5nJkaCa70Bsdfbs/b1S1CUKJXYgsR/3QvaHd5rZ/Wz82PWJG4ZBa38
diFA1u6sdtpHnl8Ck3hgxNGZaXpPzgSzY632tVbAj0gfpGDd0FPf/DeYFA3ztiYuw6R+KRIvBoq4
KftCC0EEc4pTENWBpJ6X9nSSUJIWoq0M91lnGsepkS1jNhwSmopG9OfPjyQpJefqtXvhsGdaDoUd
Re5s5H4qeNeelRbnVw1omZD9LT+E1xVyW10MWQVSZgHn18dvaJxTaFgd/K+gCcd7dxrVDbvX8FB0
xrohtoQAcBIwmVT+8iF/AZr9I3VQYwKTtmGpU2VY9nCb8Af1pnzxN1Io7PAd7m006X38tDOIMFJv
m79ZTMWBTbj93/4KbwUw0RMv57gt3mv1DPNOoN5bJI1/CalCzc+AixFdCcrICA0yGys6uRj4Em9+
3B2Ja/7iGFXO0M/fV17n7J0n2IhWZJKax6+OLasSkjVVH8lU/DlttsgbGpms9P9YeOda7qA5VvRT
ORA7/a+k0W80BbpwUtTdO/9Dkcj1JQsIDW6eHhGe7erkC7KqEQ3ZaFSqB+aRmRbVhaoHuybsp004
far/UNHwbIptdcdaE+CSX2HlYy8F9KHg9J08rbNztgvjlWge1XjXke9Nwms2r2ZGwMl0b1GAdW1h
tMjB0tmMoysnY8+f6vjK5CcMatJZsoRmbGngzZV0HZjQVHB5gG5zuVYD3ID5Ooly9Bua5vxWn1q8
Q6bCFEZvUw1EWwCKHia1GZY0smLzJN71pFcwsfO4LVSXIUGRySwpwtIt20pGhBNXsKttaBcfzirV
cUmIHkl6jDa8vhV15ibziEWv0KNM96mPb4D4U/MyF3xy2ezEf+rrDmjS2RfmeSVLOCwk8oHpCMmV
fhjf15laVxDqEHBUO5PcmZhnkqRKFvkhgXLX/Yhw2kDaJShRgSjVe7KqZiAlfln5DdqidEpSCkxh
2y1SAJeWeuW4UCLdAv76BTgrTPiuLFAtuYTZPc6AtV0vryhNTY43dIezGGTRFbbPcO7mrys8zWK5
oZ3G3/kkjyVbDjlTRWngvOty0B4v3AaCieyTor8BkSd5wOWBHLkCMXF7f4XG829rSn+fhLyWdhxv
vzVA9gwY+BiwatnN1x3QaAJ4nxpLvf8vayqkVYPwqME7yEbaJUpvqeXKGNvS6MMi/PBgQONYVoD8
7rkdoFEVFBqkNG5WENv42iMTWtHAz505Cav6ftyvwTx/GsfS8NPojZo8yHp9awZVadb2F9Wrp4JN
ARp+VvmisSHt0snZ055nfQ2AGiOU48LZWpCG0Fc6kTbNJGEMAG9oT91f1sKkueV//SncGsX56R4Z
4Qlqp8krl6agrjkVWnskrkfsnKSFQ38xyv4T1Awxl/P36bxiX8eQqmXJ6ws7KTXqOqEY82HaB9yD
+PMimoMy4ZwUwpq3sHBp8XeRPfCU6jGHbGybs/L5rn0ahHwibW5AAzQ4CAgxXbgJej2dOS+QqBly
aTiALk9w9Z4EvyeZYiDDUGhBugqFhBNmp07EKJQjm+QNQXG24asheVLsrTjhtW0Etm7TWKzvFVsu
zIDq4mCPpSu5YKzyj8A5Yt3kHNQ1JjXn+tqGSNYS0TKUIk2Hm1Q7Bh/OToUz/R8viH3fua3D38yP
Jz35V/myle/vYe+7f/Qbj4irEZ9t7ZRYnlefevUXhpIVzrV44Hw7kGEu+4+lf1ExlowroNQGBE8X
dolcQ3VQr6xbhPocYJCxlFlkBANDb7FQwxEpTCIbhYkGwTs3rCBcxtFN1W0TZquSzzlxg2bATOLx
gZDGRoBHgSJy4eCIpQfqgeAtPuniAL1+BVWynZxJNONiK4O623gLUk0HnNs2j8EY8nuo9CCCFlpZ
xk7/M9QisHVmN5GYQjNW3BhJ1QYIA2mcPRsbZ1jRWVZfqiCqZ8Jk6sH6+v29M2aOfu9Hoi+jVuXL
vUYe4hsOPHwx5yejuvKYL5esU95Wi3BSSxGEw3/EzueCkoMnUxosHraYbEoyuuayENX4RoTBeMSk
RUaQ2g0S2AXPRXjTfd1dWoDPDKo5QRaps0afKQBgaB4lul92mU8JYr5V2zyetcoVOzW1BrJ11Svb
CuJ9v5LkzF96xNoLTcLrRLEGXRFSJ9d47drqZ/c/74TOQPUeTPQDJgIwLSApAtppVRBc55+uq6Z3
nYdq/1OJ7FBj1BhDKM+a6bDx21sPXInmKmUACsuN5IIjLSKbvfiMjCBIv+G89kYn62MJ/2bIhj4g
R/KvToG+bya/UcfETaO28CllsMBTWfxbYEAk9K5Cg7wqffpfpNNj/fmda1TwX4LPvWhv5a84UGBw
htPqg4bUJ7hzlb5CTaAYs2KagcDBJTMYL03xGAn3PkxN4F0e5rlrc98aLdPWHJ6d9wF8aS9KcNrT
rQWCbnfbtqfuIWe45WSmk9qjQWleRRVf+F0X+hLtMSIBF/m4Bqn0CLaktCCseNSgfI5EK7UtBuMv
B6NujT3RRVmE1FLHqYLB4+TMcwLGtizN3XGjojebXhs1OvrU1G0oKcla0NFuRMtmSK+gUQBDRN57
r+MqU0O9jsewTXfwVnWo5cCFOtBmO7ua7Y35i87q0PNsPtnWUM6qqOr01K1RPMXxg2xPccnl4H7d
RbHsAgyLokG9WCXS4FyqMLZ/cG1tY2ZJfayXMn4LLrC1UUDSs/4UsuI+SgcmQ5i8BfCHF5DAJ+5y
2aWYpspV0fHUe/sEincQ75JWiniHa3tYc8kWEfheahhXOFjorxvYR5iXJ3ulv84xtimOjCfSkkzt
IfCguaYWvgHrBzcJBvLgcrYLBPwMJFebXQYXYKJGMsH7Mjc45Rt8ec1b6oGUxUprzc4G3Go7wLPJ
ufSEJ05eQUDBXQD5WvDnTwM6mXR2GoA4DGJAb6UEWDojLNaQ5+IHK0xLrRxLhuicxv8YyCNff315
Sk/c1I7s9gTnkDr7xFPrhU1QDGLud3whb80yWJRlkrukmDKkJGkYlYyX+VUK6hiaK6BgpqBI+YqX
w4BRWFBAgpLo932fnQkbW56GV3F5xMlK/OpmN+igiDJKxOml06YL3KiyhNydB8lH+1+iCJnlJSAZ
TsuccvTO3c2M7ijHevhZGieeUrNstcfmBkgMPcLqq+ToKPyc9bzHf6SErVXUR4aZkmJJIeqN8vk7
n/JpUa3qoKzHQNy/mBBnK2NVbXPDbtjHZ43dWSz7+4/5p1gv/+mvKmNCS2mX7m1lWLiYiqYKrsaE
Do1gCyTuF8bVgMkGD+saXHa4RxfWSetKsnPP0Hdt3mJ2sDGMWgp54gXGJhwZ+ltCicKUUZCp8O6N
vuK86dZ0Yy+FlYu0zm4mfx05MbR2iA9iiBRV69cCwYDjOnzTcVuQ/Cs1lOTF1WTJN4WcZCpFf14E
EgfWyGcdIoEoBWWm35BBDx3MwQlhyWUw0mMlt22jrD+ckIbefy6VST9yfJaoLypdzx+cpYmi3Szs
zj3XvwE5yPLcG9HdH9s9gVoVod3JqlzoErsHPfUkCHqWTiHzQSkSPKLg21ZN2LNh5f3zHIMsxT8h
PSLAsFDQ3sqUlpUhIGRHGQN//ADEToseeZ9vmy5KyW3ufLDFQNwWCwpPQdXmtpyQ1+uqcvGI5fUu
T7prAsRgwOKkSt3/Iz4+yQTpO3ZXDtltCkB1bTrxxJGLGfJJL5RotP/im71Bvu9OjJIOxQ65fAuw
BWZXRVnzPdBi7TCcgMhCss9Tc1mDE8r7LpeI1LxHWASQ/0M+UZxDrdZmZCCFXpdwDmpCyGIqgqQb
iSfbqWX+8eXMFBc16LCnXMbRA2bwVAVSMaFCnnqTw43HN5IDmiAyZVweT7Z3CRzEnG+MXyw65C5Q
sF7YiaJQQexBNjFzDrqxzZ4ip5TDy2Gyl58kPKnNiBy2b2JkeJa7V29npFzoOnwL369/t9qsJSKz
xpOdrC72RKNZG9NE/dFh+AYucsAS8e+Jf/7n2ilgGY2TLP5B2QuifcCaB5eurZdwo5QBGP8GD1rK
viRQM11hIm/8zQ4nGWKsUem5+gXvSIDKxUT/3s3ZuB0uPvDvfyrIaavi64OpNlOFCZNfjY0iUYmd
95ys1LeEEJv72rs5rFyIXvf7HNtjwVRa08JVY2FK7EVg6lsZHSwdPVixZNZZr1mBUcehyeAsN6WV
iXtO24xdDtzz2BkoWSTj6euSVUKm/QGE+EFR8/sh1uteIDZiftH8j+qlfKBKgbK8gfJH7DjeOb4R
svGOLEp/NcEwF9KXeboA/tT8DpRQ5j3/bHYOBUiWfShyFnh7vH2YWcqlpH4AbiCIOhQPe8VrreFI
9JnIYrH8uuLsx+b5miyjTgD1uNkyriQFxS8P9zpoh0buq75gFil/0C0+luPRR1cn7NxCOXVLX1FZ
4Wy84/iCqZPgymM2YNn7tbZLdxa7Xegd0a8A1kY/kqaXsRraeZ/7u/2SkSeeqGLNqDL/TVkh9nGJ
z8JrLByTn1rDqPFDHvpWhb3DQ9CkLBR0sk/tUU4otFFjQ1ZT1Tt/b4bEr509DQVB7JzWiLnv8+y1
XRuB+/8+144yM/KQqVKm1/riMChrUjJQEDJG7p6nvHudwxcqr8qpsjn/n6seUmbVz6WgRIg4ydmB
RHIQLlAD3C/aIH9Oz0nGm16nzoTR486jY7qlE9ouwkSSuMBdR1nSl0/Sncq7p7s6EGw5Q7Ku14fd
WCmcShbZflC4VnJCwmrVUqcegQfDkRXL70OK41hozhygs0dae7Vfq+qT/lqCiBkNdp60rB05ZFWp
uuU4V6qJoJEnJax15FH3kNsBd1Fb5yshj8zRYtYD4HgcO/LQmsfh31UAM8Q1x284pALuzCgrrpV7
eIetpgePymmuBRQI0H+ReLjwiZlNTW5gBHQOm+FUWe99yubV+3KR+hnp1TRqLxVinma6XYA3+ZFV
9ZuPaXD9y8TqMHnBLiqGFMJVcFsn9GdXUhtl3kxhsVr/0Mpgy/YOBT08Do7+x7Cf0Hap6Cv1dHeH
EIdfeCwHAyrMHINz3XjU+x1bvh7YauKDpyPvEPNFu+TuFFLNxmxaHsKDNkbFuVT6Z3WaBiJFKIvS
BZSK+ujZBJFit8G/hLq9I8XSGNMQahSBuY1OP2nd4ZTINKytWfFT643XVxppUrZYxOxoH0552Cfw
mwZ4x4tQNKU5eW92fclaqtKTk/eieTofgft/rZZSpfDkGVsTAksxLed9tslTWR0dWHiWLAaj0EG2
0d0k1kLitG7W4m3NcCdv4T4Xlup93r1wmmqCwrmd0fRsTy8J68SgxFUrAnd5s5zC+D0KyU+PA2rm
bVJAbBmY2EynmaIK9s2qX7u5b8Y27hf1LqpxjYmEi1DYQKYlSTfwbAKYwACZ5rrEL9OEbg9l7uoF
lyTWdOAVPZBxRSh0/Ai0xjdH+xHGxZulJqNnJBOGxVKKCSzwNDY5AuSk5/jqMqux0jP2wi2JF31p
ZYh+AuY3c/4EYY/I851MLVVDgNwfiWMvtX8YPomxiLA8g45E/O1+MOjfWd/T3lQYLL4vS7GjiW0W
Z/PXfV4YJHWD3y/VP0BGkW5LH9igdnv+UexHWcBRp1UjaeCprgY21EBCfih51l0r+9Z48UhfFXax
qxglFlWwUsCCTYN6EkQID8NoCBh/m+5dkSOd1pYqyRMkNeHoHv0GY8TOslEHLgOSqWODyY/nyVjO
h/mKGL8E4kCjMGeFJD3ZS91UuNz1Omq//h4jKVNcBZ7WcMpOkmeY54sYf/z9q63GUsSAYtUdRqBu
3HSyddl4aGfkY+bOPBw+kTux0UhRoAsMjk+JksI/TouyZMxaZxZ6Rxld++Ttt8m9NX5USUuWw0VF
DH/7pu8d4pZYjcncZIzXrdXb+TcXpsODaV+vu18UGGY5xG/qpAx3eU6aoqLeMDX93thtjz93ETOD
pzwj/CDyDJ6g0Sfdgudvq9iXxgi+ZEB40emcPVzpCdcSoaqlkuvGbFhGur3ADYKHnzWnPUmAQx1b
F299li+ac/YhpA3wrm7iPWUabW4O1VldKhtDIjTN3fyU/v4WAnouVENQfKh423orsgsiiBfslc3R
u2YgNAKv35mBqdSsKETXS4e/0aP8t2qpoig5dEwGvtj3ZWf1vIJcRLM7W1cm3eALL7wCPfZxzKeF
z5orhN/yltPQT4LbCvDkbOBaKAsmgsnvDBoklMT7Ja9/FxoD7D3909wZBUmSQtZKHhv1uDZfEGoP
0ZiHL1ylwqbzmYK+FoLhxytNyByh8UuwLFY7M0lhggygu+qGed+UFTcF1ztO/Akxq5oXnPXXjHwd
Eu/1oOrAheTSg1U8wa9MLnxrzhJQg+FXBxAPKP/038lWFPvGV4/rSSBKQRUuYv4qmPDIpvi/c1LL
TB0NkQPBkfeSBn65Zkgx8an2esQWOsKg/cR3BMEAJH4BTjkZq5AAL7mziFyhPWK1QsguzgXUGsBf
s5e+kITcVexXY/Ozp1FPUq7G2HxOkSTo/EwhVq1X+StrrvPWDrkdhpi5kHZqcYUzMuM6kqm8Z16o
EwoaC5tb0IOxhh9CBvd+ioMLy60O0oEHt1Y9OVfid3Y0481b1bxEOq6jCL/86YAmM3UXUJ2tE2NL
Xrzl3B1UXLoxRTBfWrC/0/4kEh0tlQYcn0hNYDgEXEkNbQTm631hnthMPxDJCMPoMoRZIlIn7mJF
+VCWc4Kapw6M9neQRX4XqoZfHF/McMaArQkW2/HhJhmEyJ3IbZE4IWrEdEkEb3YLCjSdJhljK38I
41MANQBrkINZEaN1+72rhQMK1SNxbdzrk9/sZStbHkIp8e57ievXJ8iZIE72mZlxrUM8v+CSWzRR
BM03UasOadp7Kbsegrow0jI3gKroHL6DrbW6No4/5HZSOCV3S9PktEYglmtLRrto6OOpv3jl1Uaa
8eGl2mykVIFzZt5aggBtQ45DThksC8gpRMDXsjW3tATkN9eTAX1ivbVkas/uAzs86WvwTdBJrJ5L
opkSUnBv2s0dqT14+8O72KYbI8GVLB+zWmEWgQrFMeLX/gIrN2JA3Jizan85gVupDiSQEnc4sUNS
f+yoDNbFv0sbPQR0waqewW1h9a2A9guAD3uWzssd/N2h70H572plLaVX+6r9a//P0yMjlJE/f3st
Jj/VqBGGYXfHFY/X6xC0bEs7uRXqYnhc9ci8AFPXakEWBAWcil+KTuQgPCODkNu1fF0VniIom/kQ
71Mea3rK8BSh9SKilLpCgAGhinLv4i8Ub5AdNPlWoCl3VivmN9l8UTwi5UnGVIgS5FFcsXLwEyXs
VZSjvMOfyEOxqJqkoWq4IUqFmVI7K1vKnIWCx+EHQSiLZQHCxjLmRUO9kL1BLk+P4thzJpDzBpLV
eDtTuMXeXX4W7fkjqM1TfpnnrFit5acJmHhuSLgdNCTiwkjNUIZPHbwmx9pnW4yOxcy/JEjyfjHq
gGPaYnKbQ5cA2hR27496xFpD9/J6bRIX5EJUue9oxaHSzUatxJ3jb18AAqzS7q0Y9GqOPpDtQIp/
fXwSlCfbN1cZHx8q7VE/5uZX4KV62CcaxfiNbKqbk1AX+0bfrK2vG028uzjjgakNm3lHxfnHHveP
XKdfzmPevCVFQUWf3RR2F+0XLO66sXkKBxKKnrW+6NhOM0iHFV8EvTxm35dBGSdcbC+MyWDJc/b8
NIoKNDAIqckSmAcGTCP0SZutMiKj9FihoKiuqKpEaWfiMDIiAn9RBQ9JpaqoAcqFHkhZY7VGL7AF
FKoyrgzFL6A9uzeCvGEAMz9ruOU8La/PN5VAi8wpyveEl4/+XjAk0ITrqfCjnq3L+NCM0Fzv3QDN
RSV4LdIXL4jcdpAmvnE7YwBDjEMHtarfo4mAuYonIZGhLhqq+Zav7bNuLZnhydFyJ6gXlKpEzkTq
EpuolMZYcYHYmuF0dmpNeAvplS0QGly/PbN13azX+kHMixvI2xRQLIyhehbL5r+51IIpxshYDUli
YMw7ipBc501bo6e6mpRsnLcOgvB0mQq+Ka40ckfzdFhFVz/IF0qWgiQ3xyCt4ngxircPsXlG/6Hd
u00Qt5kqJUr8Vu7VghkJk+wkeuCRB+L1dGeAOvpXWmrOKl2XuarUbTSpfn3N16Xf1hRWgK3HYnkx
AYx20xcoN3O9MjjWTlIXsxveQ+LoVbjRzE9BfUJqPDVrOHi+BPg/4lZaGChW0kz+0La2CSgyednM
/OqooFROJInoghLRGdghZxXjhZAOlTOpLl5TRXG1GKxm98OE1Sxq58mCUhbknfG668zRS9YQ9Yie
lQ20IeokudtwPQGMojX1nlvkVuteij57Pmd3LuO1jh7kT4aCVTQ++MSGKYu6hDGxJFzvXYUQmsdQ
MFQMmoGMO3hjIAOUBHIDPt7EDBfc3+ovBWCpWBMDQ5n5uDAhb9S8rOZTqe07UvE/4SJpbgJdCbt8
j1kmn726WRLkFsLPgeNTLDw2PljMzv5vFv1LrZQfVnu4DkMx+vVHJmhtE8nPjQQiKJP5efBpTlNE
peeY6CytorXQWRUha7RFe73+m4fWhiWLk/Xh0jq5VVYOZBnvPD0O9PJw0qJd5DHnRbzOx7jltP32
ACkpsZY3CnP/w4NafQown3uIqe04UPnQCKkEBjEVVKa0nRGhtgfgqry0qZ0yi1Ku14pmMn1Y0Zm3
HGFdxCnZMYPn6lgF68Yh/cTvVhDiqGAMIxYYsQ5fyqPn+H8NJ0OBl9nTtKPgN5wJ//3bXb+FNDbJ
sBHlyPC+P77Q6gf5HE0rCZL5AveYOGQuJKLucLWe4m34WcjQnG2lUN2qWTMDBXxE0YRKlNC+Pacd
Hsi7mp8osPXcALo7tZeKIFrEUF/MVBcxSxhQ90T2maE8L/UabECktkNfN0dz1lO1AflE39DwJ5d8
ilGqRbIpwcICKPG5f+bwvumQPOth8gUo6FxaiS/5J2AfrZommr0hJ3UtiXb7GHlusv+1m2e5rQJd
lTLWWIm9qAjR4N+50Kvda35aD45+F6smg+8dglX1aS2g/0i61N8WMDQFQESPb2aTD+HfqUUW2HRw
UXwU/zijpLGWPOspoE44a4G96CXrQosMFGtm9tvyVlpv3F+0eErsLgE6k2y+u1WRGPb5rKunsqJo
7ypQSG4DR0RXG1EXLh+oVnDa7uY7rRmHXvqwvCclIeWL37K3ZYuqKPEPPCcorLATv+pVqbiUUd16
MYLZLPWF22l+pelOtsZWfQgvxlIMYuOY1CvJa9hSxraF34XjFe1GC/SrrRefMUoVck8UTbsbqjeL
pNNyAtBeZUYCTJp0By4KKpOPFGw8q0bjuUVxEZH1oezUUSRwI/147eqon3Q2ndSupMYygQdLljwd
sw1UwDwdA3S9wEAZvazEOUloSAuzPL9bYfSHWeaydS1GZroq28X/5q6S0A09rkLdLJkDUZGlHkR0
26W/MmF+hwVvnD990aC+SFydi28ubZ9RRXg/pXhtXkijR51yPKDtcFFWxfVIYWxgTaNmbxYO9yip
lB236cZorDRl0q3th0jXAxMgqrAZRa3TY07N8nyy/U82cfnp++Yti0utFkt9lcGj/aqrMl/uzySJ
J3cbcwm2L8joTVKrIPvbXlUkZj1mJQVDTXqSdvQ64+/qvuTXOgFfTKxqp7b2C/4yq11IZA3fmwxb
yTplEyw4J1YbON7wKiY+WXGlis9W2SLfny6JHvjPOIIIkrIUWMVygtrd9T3f7pb6X0PjNPQUTWw6
3M69AyWREtPoI3/5pNkWFTT1UKTAOZRBpEA2H5hU6b0bxQ1MvudpTbMya9Zc2ha7aJoto190++PL
qSPc7J1SREHcGYPoqF6IBwKZ7vJGXVwxOg9XSry12am/81clcDKFObfd3H1bze7PVtAKQDjRcxyV
KvvSSTW5YKsOHiBUJh+ecBhIdxJAL6Qba1+TkLVUTzCU6clKOywtZuPGw7r7BCCedNZQ2oi5jV8l
HRayO5MJp8NFYyFDpFoSb68okHnWPIKYo/7+j/LI5A5wJFfnguvnhJUzFTiBhBzGxHk5zbwURk7A
KVVrgIw+NaIqRNNRPV6CKXllrSMs7gaV4n3uADhsCU/LL+nnqzPc+16nmQHe9Z3atG2WLzo65R76
mppKaRjADGCgaeGevOpmZVojtpsWVDIXQAJM4qpk+3gvwmsfBMJO0+g4/xMvtgrkwiLP3dlDuORa
NJPmAGEU3aqwGUin2cJed03dAzMPdVylAzBVIarNgu7XwpUWwutT7orYwcfdnLWwp/ID/GpU8El/
bgAbnUOrGuhbN9ZmXNDG3fyDqqJe4N+O4nlgUlZyrkI7XyryORMp9F3FYCSsyZBDgSngZ/TmORUu
oBrYMF2o16TnrYo5mCJgyWQoVAMr9KUKcEuXTFOluDxg4fmNbhpaFZbyRnKNu9DwM5uNv95OPX4j
FjotHRlSZGUBnHSmDyWSGXKkq6BZxbuHNdp5kjhEU67IZaOE2lo/W6+007swvvCFTgUJW1qS12cT
N6FK7sDz9JUqOdwyVORZkKOh/GrUXVgsYxAR+zu6hO8Kw/GuSb6bS657xzJ74+AX1IHBpheYAuFO
U5BsyW262fQQ1oVghKhoJMr/zo7PK75qZhyeacEMjzL9fpBw4Xmy/2YycPfuD4dJGTV+01voW3gG
iJ+GdpknGq64RX0QwNvUVlWnySO1rEjpy+2R31dAA6srHsMZQFMkTg5IXhd0qx5/fEV7PkNpCTmf
yz/iao/VSmj6S8U8H54huqDsIAbhj5rGRD/qlWoNNotuAZJuqRngeqjGUwaJPLjKQdvb6ISyHZa6
E8jGeWLpzTYQcuYVDZeTSSmW/OHj2xTGvtkPZiIZbWtaHpdxPmVxCrTUMXIXbPQ93D7MxQRKEXAb
A9XaBtPE9vML2GY3Y/u3paftLP3bFXBwUGwAllUkq4/e3Gr24hDhHe02Xl+YtHay6ENBaFHb311h
Mqar8Mf3/cJSsrAgo5+Ws5Lkilc5RXj7D32QkPNcJxh/OeyT5/iZOqtVm/kZ3YJgS8nO3c6VVxAk
2H1ZAp0Zrz+bVJTuBfjC6pTOJpgWrlyNz6j/uWULpZpMIan+uCPYJsDAzq8HKB2LhpjlWi9BkxOp
WdK9ypKmmrJXO2xqfldf6m6YnvircXgMwnPjrCR1DPrRrF4gT+FYDtdeSIOh++ypIZ6OKUVHv3wt
g67GHYRYQq2Vuly/rxFR0lq97JVvy+iOMIdAQw1WXCOlcEuh2FPnquHz46/PydAY7NIK6bUzlRD1
Q/syTu6WVLNrP+9sSRtgmT3fzciwsixr2j8fmEHZYsdNKmpqgIPUYeip7Nb6dp/EPXsd6lv4zckG
LhtsNjMS5qy615PYofqPRcNs5F1vuqybe3QyoNyzwUWNc4iA7MBZEtCn9D9slU3mDbP511TlHDL5
bq6FOlcuz9LBtF7WmtbsgrtHuOBifSW8Uz3NQumFn+L9tMbJp/QFvaKcRqMuNOxZfJ09hYmpYGY1
oSRUgGJ0FoCizWwGlZdvpmsZRJRlFDkUKbuFooh7iMlE3Jr9EstZcEf3kBNHfxiVDafwHnoAp2TY
PdptGSvQ8lCgq8nnj61eVXkGgplWuzaJcQYoRuvazKnK5GjGKGfEupZs5wWJBSsBql8cSYtQpMiX
wFqtxg2H8kJjTS+FW8WTaI0ngE6ICyWMrtQ0nQmh8lYzDffNsbuoy5Azv2vCiGrREYPIKjpm9va9
dqjcTKqqa2v8X0wJpW3zsMjPFQDhG3rgDaK7+itzMFA1wW9uazAaNfo4dG+jTBQteM0ROd+5Bfz6
yphvR8WHMrm5x0Nd3Mnv/X9ABnmds4df1naPlijKqNoPI7vz78G30NOKHyRQJ7mwGI8gic2zK6dT
qza6JgUh62QVkIw6/DNcLzwB893yrqP+PY7+f/g9oO5UBJ2Om+3uMp3Wa3Mv91yp0d2+GuEWyU1h
pgy15firruOpb4ODnevbU8v1SVKsCpu8DIeP+E79oz9Xa5X58eVChbaPwR3e9H2aQJ+lAw/nKek4
QvPes4Fj9ezR3yl24FJh9ejKqq6xVk2WWrQx3snh2cmKpqPTlaxIxOnreBZvnc+Feu2StciTnLNY
tup8xXskUMxufXRk/FLuL9FIMsiaE3jE0GFwYvEcqxYw7R/2ZqTX5gi76JMkceYM+e/K1OP4gMIi
UVJZ99XIGRbeqU8x1AreXURlyKyN2Uqq2LbUcl2KTez0eOmvSYBCVmIh+JyFznB9eqfmJHyU3oaA
5jmhnDqZC35Sij5Ox7PVOMTFTL/WtKk7zN5luZ4pZOYe9oLfblItBe/C0e6ygCqbyj73yIqEEB4d
XYnV5PGwM8Uncb56e4XaZ2DcdZxrqDE9eHRFFTGuTo51KjA7SGYotbhF+GjE///IbLTEf5XvEMw+
IUmlEvcsPba9Z3ZT22iFQFxsye1d/2KOMcuRyL9N15d4z0GNcOumnBDZRPZZg+0Q9zdBGASeZPe5
Os3cYnwSs/NL1MuyNylO6OuKmcjygil2d7G0DBbS6QV0nQplg1qvqImA6DMIxKjt2ZtEpp0YQov/
w+eQHdJsxTcKSTXmHTafYDAa7QlKz+VoEnPHBrI0A7QtQoXNLscoiq3XQpZb6Mjuvcfp/p1Hkk+k
GBVe13YhvqAC0asT7AswS0pkvPpgLMrAV8+HR57yp8QeB+Ppf3DnyrFdl5jVzgCVJMt9K39rpztl
NJNsTgiRRhBG1tqwKa1+RYrVCoU8uuHCZ2ulopJPvsqNwI+JUlVhIHk4B4BTs9Q6L2Lrofi+B1NG
/Up37nUUt+dH8tr/gE5kPCAURDiGlw+wwHfwFEOm1AK0tPS47J42g5G6FLu+QtYvuMmY0XE8hzEm
ilo9rLfpO2M/Jk/B9jkjVW7Ru+2DzR6SuY7gB7f6kGx8HGygO6ZhPCLW0dbggD5u15hJ+DwGgCWx
G9jJBTWiQ31JUOB+aeB3VOlLn5AgSKDiHnsaXn45LkUKmwoJTuQnjGIPVTJmou97Fzq/qxR3vdwN
i4dJT82Rjhd/7XLdNgspIgTTazHIl3E1wpFF9XNyzycVo4H+zXoWr9v2ZDVvVW3jInj7qXvE7qms
Acw9yq9GGZI4xphzqIJZa2TU03Vguw7JbHkcdulzV3hCLuUZuTjiDMFwCqvjR5vKYTyzzjWhQADH
ByL+XyXHBi/yqKJbNV+MM+xJ2IJn1RKNs7sfI4LSj+TyKTo5HyzX6VVWjouB5FNjHBgTVbpK91kh
mNai3NDhha3jGvA83rVIDVC7c5kmOBNY/4S4Sr01evGYMqd0tYvFglYZB4p5PzXns5dNCXbRvpWK
wRNAfpMKLmq6ZgoTW5HZnD8J67mXqn8BBFE7PFmPNeRyAZZ/vjQTyLbqJUgWCgRM71tztalKVzhk
IO4/nv2y9rz2CBxRaJtsftSIJKoMt5R1cyk9jenOP7527X6DO/1LBB3h6A0AhPmfGjK09n/HmFlj
ZqAyfCzj3aOMkCBd7eiXsD1k3SbGWMfe2BBZp48viGvYcrLOPq55ANJh0IagBmW6R2692quS0lHS
+4RuXQA5HWg++2dj7Ep2zmH+XJt5yxKz0OC1ULeNUfrO+Y20YpOcbErJaRcdMM0AsYjNQ9zp5g+7
FZ6sFcPlgE5dpARpgQFwafn9CVLs4q2XIKI3+atTfDyD/aN8ghzu3Jorq8KC/BrTHn9zVistijnh
+A/gZsXXw8HY259qrcl9RHp7gLSb7tj2Y4TOT5gkUKv+YYk3anfBLQ9Yodh3u7L/D/MGReXHlFep
KgZPlm4uRNIhirG2U5rtWkA6wL99qbM1Spa6sEzF/UE0GjhMfAvtYVOhrTDY1hLYj7NAqnwPK69D
SM3xzSc70AaqYAyzm6u1tAcpIJdlMcbrofslSo7LpjhDh/5lth13yODpiWI0Qc2FP2XVPUHqy4IL
E5wtYPt2KNloMmh9/JEVEcxiyCbDdYpHrEt8qr9/joEGNgGz6zP4LeGTFEuz2hUNwYhZULZcfFog
HQUvOBMgi+SZQSWZgzpF4e3lLMQUtOD4YuR3H+tvoX1ftG9XCQG+GMpFZxE9HjrUiI5bdJV9hh20
E6bBt9irsDRRYy+qMTWT9kDbsVD7f6qmq2W9ksZN7YKQCQ+4DcPRsz89Fnj03RrJx0LUICfoAfZo
TwSjGnk1pUbj0yYhcmkURCZio6UbE2RJAYuOaU9mj5qNiGPlsP88AJ55rymDs4i70IpOoWBi0EdI
eUeSMBXYACuvNk+CW6fOpVkXTYlA6Pt1Y2aYt8jsBM9xdPZxvWrLNgHV/Bcxnfz5sF76vgkbuv31
y5hQqNuZG786EJemWEMBMDPluh0WjTYAGqsla9/RjMShyhkDhlUktss+dQzIeuN67bFc+VeKTd+t
d2no+wwgTZEwXf/qa3MFgLeHGt78PbLSs8lRfPSCr345S73eJ2yt89FoDCHbCZVMf4DgYx9y9dqu
+DpemwUodIM4uCdMfAGRbQGHfPB6gSp76sCy4bnjdUsSJV5ggofEb6ObJ0Wjff+8t+Ny1pwkC4Vi
xLF4+Xs2f1LqKoey8IHFKKUi/0rJuUP9+V48Is9gjXOnXyU1XrOJ0kfMuwMX1Lbqk5Bcocqr1jzH
+V+3bM42W2LpFLhrLjiH6CFIBidC05RIte7moIIFt1olYECDXE18S8EpGvfpgdHL1DBNgbS69XF/
YH5XmV5os8opZF1+zpE94NfqoxVi+rDaa0kW4wTT/07ntxAZ87cbMG6dtjSWanpKQE5sDoFeD8lj
CPV2llvwCLRHnOgZvPXfEeuGpj7aqYJ+OUud2JcAsiEy1gs9vuNtac2LAKh4jbwYkzIXmdCdSB5I
axje5OJbd1QP/2T5KbXzY2/ErUcMY6+VHV82mQ9cSP9bxl0h7caZF2gNoIJr6RNkhUnLBYZid7lm
WEZLIUrO0Pkop0E1gUUHq/6KFKnFaXp5u4ZUZVyzZ4k7B//dkRdQgGgyqWHnWAx9TcFrSHkY5T6s
Umiv+GSiJA3O2Y8Dyvg8MyOU3/WADqvWLesIHLzikSvijTFfcQMBK+UB+aykBDj2K3Q4XlFYnNqP
lpzq1IWLD8b5TfyNJ6DlzPLLjWU5xjnvviHyjMlvG2pZDRUQSqmJh+WIXvsAfSlUu6zwsUBatO5F
0yXyG05CTM+TJGLSXdqolJ48mG1dHRv3SYegKAqYBcz/Ru5EfspFFXD+3q4yjgB0Vmmifp3xIuOd
94+nPAbXxl2Q1OBqYY1Noclit9tmjiIq4eNHp4eUznYVCM8XWi3gSdVtGCRJCt+IfVT0Qusg+rXc
KJ3s8Obzc7qFqKQNW1oGcp0NnkbxbosTXb/OfEfiwIDKiH6mrGsgwN0kcChMp7f1UWlu734MjZVK
lHynOha84dvSbyPL0RKlQUENCjhj0AP+We/98x1f62u0X8FK5yNT6ZRpjk/e37oYH9/vfBUNjuws
z7TVSA13L6rJfMoXemQF0MafG6eZHXJ2hySRrvyb0iSxyvpnktW7bOwTa3zFFvoDqBUttIJAs4tS
Q/lXpECpVP+I7LnUaj4+qarBqFbZXe49cpMQUuPVERHL7y9xP3y+m+HQDl241E/1XZQNE3K5Ma+O
Tp5dLS6qW9h1y+mBCXP573iUKNOHwZAEnAgeybDiXNo5rJzmHWUAmCY9GC967kOsLHQSAFm4Afzt
sn9xLFqsYwh5AO2fvgPzEO97SfGJnW13AFnWJisovdmGUKjH4PdrBrg1TEfVznr0tf5nDs8c3GMf
kqq/AklIagvUQ1EI5hE6wYmxI5eoSfIDSv/2058IDr9Z88PL2f6Hhz6KAp0T36OonXUy5bONX7yw
ytQnVydIHDlsSVyk8Kv/eGquNgbxYbsYlWJFNc4j7LFpp/2wqIMfuAzch86F/adgAdRLy6pZxVxZ
yHwtU2TULQ445ISI6AT+CKjXbbVK12I2pkaKO09IXJOVvUwQD3MNTsAzrwXeGcjpx72fE9m/PfIU
ae/KRr2zNA8spbPa1CTVglK9Mc7JK7NPQoayCL9VS5dOCKMYQMHTLG2TFHIpziwCemSDb9bhNhok
yOpcn9iuENXOcfi0LlLls/cv34XoGXg4yXu4EZVOuAYkfFL2UPCuBjdS7Zw5AH7gEm/wM2h37cGC
uR6KDeljM6j8e5EXJ/ji4wq10PkvD3AwoDvn19z6gmrRbUgOTcnG6NukMW2XGkm0FSbJz8h3cndw
RdvH3sqzC9apJfrA463BXD2Cu7pjrU6ORjK3nhSd/siabPhY72RUi+vZcwQJEK7NGGjZAS6cGgvs
ewDNtpZ1yvuPUJz6NGb4YFUL6ZTu7E1oi5B2ZIbtW7+RD2GVs6Qut3XWnoldFBi4bOrFFhzZp2zq
yUaMgtq97D/NhUmrBO2Sz3qMAVD8QYn8+IPh6suytyVszbcdoscz/6a0vjWpSUaZQNJWjlVB/Z6w
mlzvrOOUtZhLAmDlG0shM8bTIwcZYm/s4duI5wBED5WsDzyRmMmVXmFMnrmK35oMXXPraWWrIJPO
fhrKdoSppI7S2G9l/YTfp7Op8AR7fXAufhB2ZuYZJs5YI27VlksIFdJkgG68utGx/svAkxc2Q9Vv
JncfeEzcJYnsCmsmHwpjiifJUeeCK3FEJh/X2xdFwdh9NmCqLtdapbPPFMhNq0NJ0KsGLzU9BMgq
bm+VRyFZ8LYBTRAf0mmMW9jCu/7JgdMTOBPCQGWNyz6JgSRI/sR9fNSKrCo57zZRwLFjJP3yobkm
n/Cl5Hfa2ySPhP5we9ddWO5/lQP9KFlD7y/U+6OkXCpguEx7xwWvrht59gS8s2DkQUIOzZilL1g0
V8n9lgXBhzQifNdU0i/hJ/W72ooHhNOUXAaDSpm9hm+R92aPvIsmiQRpe8pr4/Lf2hhbyeBkK8wH
a8SIj60VTl2VGkbc89JTAMnNwJmUaxMW884Ugw+PRhO3Ghwb0B1GwgaT96FX68GVlw0yeGl7SqzG
2liZKVQ3WWDPcc9CU58HJj52++c4SWJSEiqLF/3RSOGQ/8OfevzJGshHGwNaRzQaeQYZ50KRCGC3
MInuCF7uNZhvK9uOxmzAf2QZsyNKUGMrl7rxXB+WG7n1LGqlyycwQcrLETj1JcXDtkH/TjbpGUPg
QJcuJVHhXcT1zc3SFJ/RI0mifWoFBLxMW6dCt5CaZwoxkkoGrWkVuFDuOot0TaDiCHecW+jAFqh+
d3gV2fPzCp0klYD+8ACl8pKjsMMPa0XyHvIuNbAXSP1K2SBn0mDwaf+ygyqNesEWYjVz//MQjNkN
i59HmwSVVNek75MdukvthFy2erOWaqaUpHaBNXkRRnB6wd+ClOx5eIVjp9U1vdW048DFMvkzS2+n
TeTxUBsWhoO1cOYX8DFkpT/CYBc21+JQzgvaayJw8UVagc6Em4eARcHDld2mvH4yqpy2djiztqK+
th+JS/fR3sEHWQ/Bm/pOnlHxNfE0fBNVuf0r/oonBtG4zm860FYQYniWWOIWzbHmeYQr1X1Cs8sU
guTi2/bmHAzrI0s6Cc/O5B1CWTxi1kcyVohfNP8oZOCSM6IjiQFnWgxBXpZ0vqVi8SmBdcW4NLLQ
EekDIz9534Qr0nnIFIUFpcLO3MaE2DVY/EDkAiXDC52pfvH3P2CGe74KOZSAsb8pVZyR6ttt5qGF
vGLyvd4ooWmHcC1IGhAH0jppoqoIgKngTQWi5nSWtxtdGRZc3m9ZmtnV2JevOg3Pxq9OZEfwru9d
Qk6ch3nZBdRQUKMewyt7lx6yfYam3HYQc26QfTl2d9+MHJL9l9CmduzsdtSdCIIuJhZX7RVfCTed
u7LgjTLYaehVz53GuwdRjWqCFZcsh6lLl0KJZHzUjSMyDHk+c7OMdXOCK36JpMYJ2zqq73lWd1Ln
IdGeVU3Qc9j5eX3PiEBSMro/PnQziBBTIca4YYBxvtKKPu2XqkWoA/zVQYGP9IyucZKlc3JFcguh
ZEn+b26iibqXYLGPwsrhiGuRXouQQFO0rQBA3JMFw8Q6vmLccmFm2I6Vo59Km0qpyO4QbHwfeeKx
OmR9fmJOLWnQvP/1BLxtMAobKW+jQbSEgxXdjloZUR0OOy6XmYjkyK8gXMSKvMgPqpWlENXo1zgY
RU1CUPk0U9zixLuhz9VyB4+Ezfv/8DkQP31kMD7n9cUIh9j3YYQo0gzTiBf0Fv1pLvZBXPgH7ygq
/AdagD3keqUiTKY9U210HrQbtZRvZNnqfswMtgYL0KkjuuDfs2MOpZCNOQff5tybs5QHrIFxSP2l
T1bLNgkKLwO6k+H2BAUNGwWhongFQZf1KwTOqXE5SC03dtReMNWqDdCkaXI4oJZw6jSUJi7gCqXN
AdPz95ieEKDmPnROr81xPXkSz/0fuK1vDIYr8ppDQFxKpgJwcpFIVqzXoweLA91sNq0zZJGX3V+p
Hh8rAB1bhsg9YXnC/AspG7KsqxjTCCqH27fsJeGSPiaJdUlHRdoK9ac5Bfy+VDy/0OrcCzSygd4n
fmez8sLSKtrQAI0EJGf10OhGPXmNIi9oHAz/XuGt2lY0kRtY3+bGB2YZcaZ6kfoOSvs9+9eQjrtj
i3yybilSzKHoj8dhpiHfVXyTopbLwFZWzL1Md3WSW40kElbDf8ooiTK697LwfpnFc/2GkTBh5l0O
sGLNee4OncyqDcZSfzNIa/YFvLJopKX9QVnU0dru7N2qUU+07sjJFJDxqg17N2LZmJuAx4VdHb9v
ERGwMMymjPQH1vBZ/lvYCVAPji80r5pEbLs0ML7aDMXObBwHMEO+p3KQBI4Rh2mTBnDAE8EGLVxu
YuaUNe1K7AepWiNx3WOZAL6SRv6zsdfuP6LbfoliCqrjEfjV7TTExT/hn7TRM6whfSiHxmzx5pnI
rMkv+I4xEm2AyZqJ1yO70Xds7aPx0zxl5GldHCTIsrSsSSdGm1DkrowhZm9NTniMNlIyYtWOhNxh
sDUJq+cp9b0hG3uCPHcA/rR5k13fKOqZyT4gpGvhCpCcucoOuixGhDHML6Px65D7WCZRTTFMR89L
2sOzVX6s8Zsa2JwDNUSXAvJQO3zBI/gRYB+Uq96XyC2PVMcB1iym/RGTFuZSQqMNUOik9hEVT+gi
4tAiR5ARA/L4UMmfd5YN4nK3yA43A1B4O2aMwbVb7urdLi9hSP1CQTHXGQtIUQcLWqOgec9pKLdp
rvUDX1svWv8q3+CR0JYX+VadU0FZTdV/2/N92oB157kIB+xba+zoZIvD/cAiVE2ISh02FsqjfVpB
xKVMhhEEoE5eDPBY/FZdrvjCQNdySB74A0rbrHlkdllokmdZFVGZgLvFjri6iMtQovgLS2cMcGEV
o8sxMPPmgFJtsU6kthk3fXsrWBjjUIIzJtxedVOO0sl9SX88ELHNqblkFvW3HTPG0l80WEiop3yy
yzPNva2PGPM6ArliS5A1Ya+8t/j1fsK1yQNNmu5pwNaAz6smDgWzxd7BrVT0MTYuFrYzEP4FI0Xe
I8rbOsIFJv7jo/GmaZwN3Tf0g5jzZAHL+biZT8DyW/aBqOYNwvHs0e2YxK8rJ5QCA39PE4D/VGRs
qCVBv9xCNvizfVUdfPxJJFGt89/k4Wi65GK0LDOAB9Pbhv3PNkR+ydsqppazexnJ2kKvRn+a3YAl
45VR+iBDBAydPNl9C83892+C4cp8CVHvzX+QtXZdSCiqVXcDq/ZGFMHtEKOIhz68h/rsarHomQvc
sFli52ov2nqL7L9UQENKBQd5VJ5C/RJGv5jwizdiWEA01ISXMg69zve2d5aYQi7mw+WmugCB9prp
GF00dyHCEUgiO+pFw2oVZaBxPDnrPLybr2liwMYXZsMQSUYHJavrKaOsSP93oXbdorJKTzc+pKT7
LXp/L5+QR/pcu2n5HYpxHZjUUhbi/AqRR664otP9+M9FGdQTZPaIrCI0pQicWMi0LE/XJTY65L0C
LjtcOdD+cub5GFt9d+LoAef/8kI7v1/7ONRZdW/MdD9hwcty81NuDyB+f9yZATkWJkrAfndCpNsR
x/mIJ4bFY9eSPeheqA3ILdlSm0eqkfIv2CgN+X+MMBPu6F49WUZNU5xUR5QtSCaNyvwGkT9iBuqh
NOeNOnmWFOAVam850n3+QQS+gBIVkSfURzPAnvZqQkCAvJaxD/lgD4o465qVAJ2rGk7YwUd1YNZ1
5PjyPOjJMO4re/vBDvtw6bCZsXI9I+0YEH/YZYyDYiBYzfgquAbMfyTUOqthL/fINJc5s2WnT4Aq
5+eVhi7rwvbI5jrED1P+tUcSDDzlvFPuDgepkviePguQdbNd7MdhWglXqzdEPM0n8VovAc5hw80r
cCPfmuY4MtVmviA1DJZH3zzDBzKa2GfpcZqhH9YXwi20M2eWIpRjQivVh76nuX8KksfQHGcfoNdx
1gec9HI6dPNBimjWOK5uoe7qH4t5+sK+xgJ0qQv9rwYqUDChiIzGipNoztg0WamtvuZRMoPwNp7p
tLMZeLd7e6myDLmyC0pyy+IoHawKh1ryWx2qtF+mhOlysrnkuiGIjsX/x7TUsuWMU3OT/0+O01Po
U4dICXZYteFpLzdCgVkU6v+JW87GTVBBvoKKu3X1NAJ45NBetdHRrkFVEVLQJ09T3e/+AndzdAJv
sdNwO6ExdHKWaJH8Oxwfol6foYnyTQ39A9UeLXDaMdU8md3wl6dW+jdHFhkbQJnIqGARzR8ND5Zh
tJgJj+sgjcXWZVPMMH+fZEsdxpg7uDe7GYpxDDcTCggZf54A/OsFm40gvJ9eQnL6tX3gALA2kgq7
O71LK67GBIAXnAUsVdc2flNaeIIXCgCtxGikZLWNTjrrAkYbI8Nl8tjM0/qdjAE2If/EdC8TpKuw
cHME96exuORdc7LLjteSRLKK+eiZiBmLhdBCwFVKq5TVKGvdyHZ64Ef5+eXU2vjrbDdfMafGlVD/
RTu65lVm5NzL2abj901s1KRMGW3+lMwCFLlDICN1FqvgGq4+FCl/FMtSa+AasVX+6ZnfJpPEqVyK
n1eQWFww4f8VSdo0irKpjGLy9KrYWvzpbDxU8a9UE7EfDn5HC4y3bycncJl0+f8bjrhemnFEtmoq
ftP/tV2uq74cy1AGTMeY01fHS8jxx8mS2Qb6sFRCpFj+BeSDuhgMAxYXO9A/qICEIF53s42ZtBvt
iCdJmRO/9is6Th5IxaN8C8nZUB+62KoUQjOVwe/AlnFdGVf2YjsgosMpF1I4sEx5G9DayO6BLDgJ
digw6B3WCetpPuoouc23Y9eBkJA0fXM84k8aiZRCGpaZfytDtq1uSIWXKlbh8PRgG1YoI/nP8wZ0
pwZDviCFW/8jQiZmMTLlzK0bs56FCD/QCZ9y9lFbS9nRXuTVTt7ppQU9ZyfgkhtQ39Y3nwL8tex/
Sgmuf5F4Xcr7C7uQhzY2FQ1o1LG6G5DouAoOSSr+vFc6iwMOVJjTK4awhj+s9CKw3YJYjQy0CKAJ
hkGeoI4iCBJKsWVPabqc8ryI9+GDgJhLBpWggI97zDrJ2zSrkpOYfBEgDlePUG0icDieOH21jaSD
OZGhFQ4LXfSXshqqXyjojC2Ee2Q9w7yMIFoF5kohwkX2hHBhJZkNszx3Qx77qO4SrBX3wYnAU6td
YnhLwlVuIQG4O1yyzgxZI5RebcUZkxti+kwLobKY36n+0a7St7vXWOSX/HIcKDJf1+IJhUdiCLm1
YPRRHZ8h1U3A2V2BrlZADZ8CWR0+yXISb5nM1AO1XNN5+uxpObzoakMsSI7sUAGqViy0KHhDc/CS
7J1N1Gh8PYps+I1lKeQonA7n8VC75gNPAu1CU1UVc1FPqmWbo4HxG7gkaEAydOBowtLTA89AmWF+
un5b3okXOL+Lx1SS9FE98dt9iSDjhBczEGG6eYwarc7rNYtIv+vydZ7zZk+9YSxt0duKVDDVHijp
ScAsG3ZALA2bhRccIr1qmLiEgUEmKDHQcvb+KCcAPt4xl0Hs/vtDB/qsQ3+r6E/TsJkd/0NLe7cr
b73QWWQNPFI30mtK1iO+VCal3HcR6EKVN1rYWbH9RTlVwuoQd9ImPod+BktsqsrN/wnLrwwHx8p1
zDFn/tek0gwcDehXwF4S0yxcfQ3rIOC5IfGdgAbvQYRLV6bQJFqCrqHYwPKj3PWYQ0N/bLvW+E8b
y75EKZkRwY4dNSOo9ky8zGelbcO9WizUWkKhaqSRcXbTjhEi+w0WzFJA6R2CV3ugj9ie2p9/i49E
aRm2ND64fDexfnojJ3ijWRP33mXA4dH3b4GtB8dwUNP/GXLacDFCqoCJEixK9lSF0Zt6gtNeDijU
D+BK5rWTl6h1hjpj0QMglSsxwwkLXUdlcTjwcfeko1FfMHbp4LhSJGbkVdxxuai/ZAhNK6huRl0n
d9cnaQb8jnMAYa2+ZAiWAzzFyY3PmAPUvIRgNHw3BGhc7mGLgu9ejyqx8ObH2L2yY/Coq+XXXSro
iwOxvDT5rQMnNDEyOVgG5Yy41Y8Z51c1PcPOuXWQphlD0gMwIkRPmmpEKQCJe2IQjAUgae9aSFrZ
hQ8fkN9aRfN2ovMAK1e3Al2BixS1aRPByghZKQhzvqyVukngKiarg0zqItxzO7IvbJv5f3++HueI
E7D/rFu8sAtcVbzIOaauRO9fqRSzRggoAkBIJBDN+Xki0AXj59F9LX2VmJGr8w0aP1/ugv2oK6yQ
PnZzbTQUdygodmx6yWKOK5mcjY5jaWtOWRbBFTm8of7ysHeCFjEg8MULaBTY0uHALQ1uvNL6HQlX
V9+cuw37W3i15wsG4c7B9cnTG/go036CgL23V3yAuJ14sumkV4zA1LRjgoqLaDMufIxqV38fMBKn
rJBu+ylVVrAMm/MOG0m/53PrcUGFcZqfXJwFyOVXLML3sSmEChb8XZPLlRnPKwmBx+gGADHFPwDl
MS7ZV3R1S5j4sBh0kS9MR7ufGVxMc+/vVehxnXqegMw4Q7it80GNODiQlskH4jivySrPM0200yzw
HvuoyGCTPy+s+GmPKtrjJWIvQ/z6QA4jzV8DkYk9Dhfwg6pbAfRsfQoHu821k22uBhU+u5tO+sZl
/YOXUfag1WBsXdh3oSBtUdWHXVMJz5Jk0Xlj8Pz78Kwr0kjv7bJatPkq/KMOsZM3jNeuOI614Efx
nfkpepEWZ2k605NgBw1kGjFLZc5TSatywOnVrJ7VgumkKk01+HRnojISZDsr0GiAoKCEIC1h93kF
RKSLlis6gp9t8ZNiI54MIE1Ww9/Ht/5pLye6IoRHovaSkGQf+cQhuiZBzoUY3wpZFSZ5H5wJfhzr
vNCTPWJm/MtzSJ95i5GFAp5AwOCtKXyEdLHJK1EVnE8f+/SqkCRvxQj5Tc70e1Uzepzhbu91iA5Q
9ZKsdsV4vjdcGmQHkf1u8TldXE1NGwEui1crIZ25hhb/yhmMsQxXDZPsIj6JxnNlpHynaXRzxpB8
qivUbm88RD8y400C5ZG/xzwLJxylXrdCdCVUucBzf37ySjWEUtY+IZY9qZon9v+IWrpRHAUiZ9U8
S4NpQ+HHLbB+2xstxuHPSLGjtTOksupeEGyeEyaT1vzazP4DrfXJgeGvCyTKm++1npcdWyph7vhf
I6CRAF5ADd4uDMCR3Fk/DTsknWmsIeb3SvyT1+9Hi2hQ6cP3tUMuFTFIuzKPHQOob19c0oyDoWga
rt8Hw8LyD+dhs9kMIahkWUqUgkTOkN3AOHK8wXvjPCGMMDOsbZeuLxSNa+rJg57q0z2ggzo6wN/E
oO7oDHllO5dmT9fk6QyiMvBh6ZH9V6n2XwR3Uqlhft5sovT87uO11JxaVOBb+m6iF5DB+QqB68y9
mrqbhKhSvB3fv3ykhxcZV2AipiQxHOjyGJCsxRrlM5ne2eJ9d6C5Rl82uECo2y333g85q0ukh0Wr
FdbkKtGEHjSB8emRwePQzpD5hv9FU12H6q7uIOxnQfJmTjZb1Ubo2f/k1ne+ELtzrssvMKsVewxp
698dDtkesIMbKqXEwLVH8XFwwzUSydfLqQZwcNPt2MrbTL0ySnkNZWw2nhid+OPef6p7C8ciRQ0Z
XlVOeb/rN6fUhrlotzjhpn/NUCucEzaXenLZwyVDJMLM6EDkw5yYBbiIVZR+al3pIsgueQRS8N5U
9mN4Wt7s4ZcW0sgbJPN5sNeB16Q05sVaGK2+xmfYvo0dwFdS2o9lFxTRvPoQJRLD0EjqFSB9aU2A
YkIh6Sj2LKNt0encVsKiovS1/KgAuA/d0NLS6me6+2neOAkKYZoLsA38mdRsouoQPZEMSFLhJg8G
+o46VOPdcTxX8WweQ5rC+D4cupId5TmWq48cn4Fc25e5KC2KLiCNd0o3BQTB/Yy6fhn+GdPHYOKq
2cBqJzJoka8SmX7wBFyv2KiXMcivR2vgDDySE68Cz9UcaFOmxK+aGqG834yssx94XMEbWoM/S6Ob
vD1bDEy1y+r5iTLok+ZoIwVvwGqxUhN54l76Xda+mLtnN3fhgaXlCV0M9GLc1364ysLfo3sEG2HV
+z+GRUhK5t3WpcYoVsLt39YDFIgqu6JgCgvUF1LDjy7iYUCAj89XqlRbvPrWMZf8gV++G2FMt7do
/rzZWqqnjou9d50UywQ3fMqfaL6rELA0pf/yrYlrlZWTx2glikJCHwMyGgREFdlRIYQhuVkIJE9r
GNQqlr52fBOGSyUhuCCcBK5bkOpZ4LhMCGf67cvvJU4YA35s6Rx39OyPBsAznx5UAHjlq85hOrSf
tVl9FMEbW4Y5BtleKr1NmUw/cQoK8IWuElXgndLwJBlAyO962kOGj5qMuOJwNfAjYItrbopa5O2j
xk82V19xOZ8cgB0SEJQzvRHMzIelrpHOrTBO3yU0TH7/P4T9l5LN+TEwqueWsv9oW+x8d7XB6O0s
toxB3E7WpXyutCYpVXoRSIIiDgecdWgvLL/L59043W2lGWtzs3LgAJIVxJJAOnenOpigJ2QPr9Zj
DHWBIW4GDYunQnich5e8ZPKvTnazVfIQt066JK+iYlEACgKW3BXcTA7hW/COxxGjlOevo0w3glho
zh8eUC3PzV/NN3yxlGgJVJatSWg3CWX6gAmomcPSdTlGoE7Re8G/F0LkMKVIXGa60OP9OxdZU+Z1
7LJOWz7vxRiMfH6PpDA0NhqZSJkeMSFKo5udzEWxEznX/05TJKeDInty5CB01RbjyYitcnZYN8Y1
+Qzzrsc/nt8oCAO6twLhROH8I5XMLCt8hk8MgdYBUtYOX/WFQjLmrGb+b3tnrXN8E5ziCPwdTXTj
HM19MXFId1lE2wPO6ek4Lys10BzB9LeZC/LEzBo0sfu4N3up2SZhLnkSmj/VetQUVKtyAOu+QCat
KSS9mmiBb5f6Pg0ESRt2gPYLlQU01jo4STYB/D51muSRXdWcjnRunMH1y+jC4yEFv9Gq7gcT0mp7
Dcv5OWher/bE9FOAmTQ6MRG6HNTA4NmmdJ5GGBClo0G81OveEzcIu2tDLjBpIN5ObKErQVR36EPy
LMSFFlAfKONnnRbRtxMDwdx7qs3R5d2BtQpdk9jZ5hX7fZg9BTurXKSnJrG0skQjX5SJXMOKMsct
q/E/fORo9JQowaNv9c+gAOUdLRfd2v+aCF5ZxO8/oNnhUkhmZfgAz6Ht2yhICr6S1K5aASuI8M7j
EfuAWp1c3tmfhopUjCnce5jOTtgFjHp70Q3znE6cmQXxBqwYLcuq0Ln8DaFFv5SiOkKVoxakHS6k
876GEZkYzh59p9IYzzIB+qmuNWHnhjzOEx0HsRdA8sgA0xhtUHpb5uASvhQm86f2aL6RhQlhlv9I
smGP75+G2N3vyYL+rzWlpTztRlFr1fp7Cl/MkWB7UNGMXf7nfVkskSBzcZ3OjJoRO4bPBm+LRTzR
I451oRe0e4BmPqqdKXy50vtKBs+5rbpsKSOF82l9AsWAGVBjXDi/vFFrc4xyc2oFj7Bs2R9CviTS
Z2vZxRBLovT2NZa4zqiUnimjFMMAyFmCtCW2Tp+G/lnNk3oiw5yzBIzyF5GjYiR7DEY3R9Vjrw8E
ee6VvHBins5ORTPDC624kprcRpmk/j0ebYr9Jw8q+KaOUhrxolazn2/QIUfrWfpx34LRQKEuBKqR
sD9/pMI5AUlLemlVxb7OQVGhsz/E1RdxgOFvD942CAAPesEVoPkDqTkGjfWrI372irAybOSqxuz4
cwHAc9TF9ht2OzVXQTeHmPP4TfnFM/Qa7CjxF2v3AVSH7B7cdMMVfR6SrgnBQLoHiuD8T9Nq6qGp
shhMNbNzyPgxmkUxABvzoPxGe/dY9S4/1DtBnGqhmb6hY54BNe89Dfw2e8Zkr7a8/M7jqJk0gDps
P5cFKkiYs3dhqOss5/mu3/mdHl7TNhfMDGKP0rriAM0iaAMW2jDI9dQ+gTDVyJblwPbMcFcUwyxZ
GuNdcChHh5UXptmP6QJBC5vXfKSDarKc1+6r96b9lT/RgLlYElcEnAp1JK4s7M9HDJI+XaR6Vcet
wdrB5rpmT1ycishGDf3sYQ9uPLFeIIBuYY1+9hSbtUKdp1CaGH6imyPR0D/d+lqbGyMo3UEzpQSd
4tkeFdfp2AgwSV9FZOxVzh1w7+lxSH9VJvNhXwh3pRU1wnMiC+lUIm66eIXKC09johCATehdRfcJ
GztXxZxOxSXRpqBBrUIQXy9h52FOFCJzmtygu4+SXUxLKgv1BEs0BMHnvMGxgiVg3RcyuLXKpB7S
4Zy3pi+6AXvRDfDRXOd+41VdQ306wrn8djz56iBsPN9s3ygq74dodr2TmXlfgA79qX/uiisrp+mI
w+MLXq5KxE5WbG1hh21kgUAkOhTlfr2G0oN8ZH2YSVekaUvnXZosGxamMDCkYmx4uKb7LwnvIjiu
Rm0ymdiKk/v/DBh0sWstLcFHHDp3aYkThA7VG5CUgo2N8tlXbFtl6NP85pCvwX+a0SO0/MoJbvA9
IthQDPXHu1XWXmP5ySojhuRMaDDqOE7q+4xFuGa+2JmScPfL7fQkfDEEJizpzkUfU0mmBnrB4QpM
5F8pXoJZcL4Bz6YwVJGKlBYDDjaH7J6H2vhSFYxUdDrByOLqry/kCeqTlPI5vjaZqPNk6uZ1ic4t
zn30JcpMcLMPd3K6DeyaP23ae7cysBTwHuAbtGyahl6oEdPOGwitQ+azA05Sb3BiTV6ZMAoGr8fV
I6E+/T13eJ86u6QEzuzERDkHkhAUx26UsYnRvEbmW55LJiig5jJA64YeSz0k86nuCB3WRbViRkKM
VrKXja/o8s8r6IFEvVWNmPiJrOrgp22uUXdF0bPoxuACWhe96xAwhly57jLDCsrHyyErTnlZa0uI
LsovUmRqGHOOZynmyWa4idOKLrX2sni3Qw8zM+w2EkleOK8t0EDB+NH3AcitAnrYR3Ldj9CTF6Z2
P1Z/LLYAbbfYWVLKmyAoSnBW39pvno/MjhF0Mry6f8N6rUQ3dHRvhYdRvNBDfSnaQlNfViDTn7VD
V8sEG1FLh6b0afqyk8mx/0G/nJ3zahXiMwHSnunsaYtDugwSMPQdJ6680821vCANcvJI6zs7/S7t
dmrSJDxq4Ft5BNRNKooCcTgy/ongOLIxmV+0oHKnwLpwJvlpcUuvp1YkvVnVCVa+U2mJcaxv84iX
zK8tH1euGQ40flInmqyMh1IlAUtiwL2y4fMb2bF8766zUZYXmwGtLAGh2Z94ixNdiG7m3nQClHwn
D9h2sdQO1cfIE4iJhFNH4gnwDDSkC4NskbSQN58w+sfoRVvbsdfMWcoH000x81kTYOJJikywMRbZ
NpteEjFybfaSX7FvlRV3T8CZ6KvOKdCGtFdHTJ1A94ekT/yqeAm4Ww/8TFTKuGcwK+YKarGte1dG
HvBc0M3ry/EtWcpRHGCZRr/kHoa6TZq+Uy48EiY5hAaFkljRmSk10C9lw8UrCgInKZpjYPWnBhoM
eDDmQn231IwBuCsF8cIEIOMuTUf7bhP9w8URog9pRixGzfYcLhpBU+0LkrZc3jBZoByQGxIhdLzl
sLDImkEON1qURrdXGhVXFuqB22rCw498OKrJgy/yqf19RRLsw8TCGqyOuQGXjy/DLeuXdlRdpyt0
1v7VnI4B0O3nsg5BsSG97qVC+U90byPho1D0xssylSFE+qpcm5vZhgVaOapzTDyqPKDDxfF98WZl
64slEgWGXvghHdgCOfO2F8C4sb00ZtIvvWaHZJWI5SjZS5mEw1+8hrMzQFsrpecv0vTOWnEdNmhU
Y4kDQOrbAwNPNrWueEs2Nj7YUqbkqrwUajn4ggOMfv2SzMGO+YLLBMkTgQ14ALpPx+gnv3HeMtqW
UJi4kLfawJ1e870xm01/KzFvpq7gBRJ2ThDg5Rdm6LCico+L/wPw57o+LIjvPhYSVVfjqbT6uAl7
ujE4sGSc+B5abX0m28uGgm+rAym76W7Ey0YCq7KaHQxNu3Q1pCVvzQV8aiQ8DO6oqBsXa4fifbkc
MOpGHUyV4KtNlmAKpi5JrvQAMalHEnq7gS2hCkLr2Ns8Tn8xd7GuPTcYaSfN3E2mhIG0XQe0OVUl
95ES3r8Y11VX0e0H15KAW2ZUnEkU8kywJGK7UV09j9botnIwqIO6E/APBJhMUN2QJjDDQ/IyYu/s
cq3kn3ASOzJAH67wK3R02//xtJMiXGptOUvSTMHwXeVv6nBMeggJgNJ57MDiP13oUl3glNqH0B7r
Fcc4WPq/NwFh46zYPvrPd6SXS+nH54DEShmi9TM9UQwBNZccaEnQH++rvKB0UvyyUqlyXWWVDGzy
WBQmTBqcENRYb2K/1TStymh+51fcv/+tEIUMiC6aPxYalB+qR/3B+5okpfvrYGn7ix2+kAc4DoMW
fFZibc/kWvRZtj5FpLtZTCst3BztrwFGJkaFQyZaGYVv47NsKAQ42yIYkIucdGfCWUS8pqULYUBL
VtlkysIs7a1VQL2jMMRTt09q1OlfPgkZ067x8KtTIPKRye7IcgrqJHmiPg4NVAqUUezy9sgmOAyD
3kZ6M8FtSGBOBe72JAqt8rtEHsTH3dSRS+xKfuhW9qgoTIqBs9WmjuQJEo5vv97vv2FB9HRLbL3y
sszwtHG4wTTzfsq4YnuWcA89239ub101DpR17vEPdcJ/c8fn9JWRjOmLwBHrdJofUIFThzhKJzyy
GEtrNCWsaWqR/Mj4bow/uq11y5yYWVmozy5hqoX0AY5fRnzYB+2Sgzx1nCPobjuNnV9QIwQIsaUG
Asbbdd9A3jhBeyy2jKONq7wtE5/g5Y2WSAnFSyh/WU7PZ8TCZ4Wo3bjMgO3ChIzh8aKtgXu0oza/
yIZJ9C4ypSibhglOxpecazTJIUdv+rTIalMCpPpTuNV7dBRSQZXpMkoc+UKa0/w9BRtHG1PEQMxa
eTJuEuVa98dm1pzGw9DcrNeV42QyU0WfWIff8z8ymPT26jkBEAp0Laczp0gy02mI+NDDfOOVWxH1
V/JRdODBRoNrVnna6H+bM4mhcZyUJRbdsKWOAdif4G5+0Q5fB4TtcMKiIIlPPRUULEkWsppZQoVP
Iy5Cf0lHVBVYSGvKjwgam9uTnPqUBKuaQ/h/uTsSUFn7f6q6yUSeZDgNLC+SBlUO/Px8XIMCgutA
O1noCytfEJcKuw6MtUxDQi3P5/N/pSG3WzuYmXTRDQUPa307+p2LbNOt+MK2Hx0A3RLUBwGqaJBY
R6Aq1SKRe0qA0aqAGY2hdvbtrLIDMyQfxA7ZRGS0aIhrZy+8SNlKd1m+nYLxCg+jzyYRz4TrNigw
TS7PYgdxoVQPOz6SFrkIGxioOSFIEPMHppFYzyZw1BX8BcIfcI5E+rtOYmobG8n7tze/PbD/q6Zx
t/m3idgBjErfYXyBm3/sz4VxQuEgsvnZz8SS5ZUJgHZ+0edB99o7+5/aLnAqNQrJTAk4xvk+t41B
reul2XVcplcm6Y+V41V3hFpmkW9tchLVl+Ar72//8OjnqEktasstWLRS2BA1PF6c80ZwPWkbEZ3r
V0GMRT6EWJNxKJ+LRF+QXKcsDjRBojJuNSFF5lp6GOyOrRElPZ2syzReSeYIQy5mt3VMvpHI3UOH
a7zek0SoP3Kv7dA5GyX9IiFpuDaktvaBvUVh5bNOUy0bYDTCB/NAZM/Bj4MAVX5vLNsC3b6789FW
xcMHaLdVHLGBMWwYJrQPvQOzMyJqbCV3+8dCcQKEOZ59xYhICKDkQdgjEvxZ0TJG+08vaeoNA8yW
gGZAjhwzdZl2OJFAeQbQoBg1O87LRw6UrL9cmxTS8TQmZJfF/XI8eCb71GC/EnMHowyEENLUOoE2
OclPNo0VDoysLj2XxT17IrXXD4Dr/oB/PFrXXuM3HHYJ841isl1euQQ47M21jkP7wBcN1pg3DzT9
4FfbLV6W3iWJdWgpKnTqT5Apd4UOS6hJcDeAURXRzuGNjU1AQgiZCGA2R4/rxZvDH3Gm5suI+wTK
RMsnBRngXfWSlbBoLE3wppRIo5o3I1qwUy06P5G/4M8XBJ8kdl5BdfbxcTP87EievmPS3HVMDex9
zxssoKg45/MLYgk24aFfpGgswa9aAILeA6DVmSftoXNunFLdUWGlDLE5fmfyIPHZ4DgrRiphEMv+
EHjS2wFhLRHHuJUVKTnj1hO9loE1DXQDt22fvEVjBq7yoKHVtGDIFTI0fsnNUxPm69X27TI/mVxu
vg3wtvaQNv8bQU0fMliab+JKrhqDsbWtArMgEAdvz/ZzY2y1TViwvmJ4aE/8i/1oPLdfi7xXzmA+
FtxAyfiTQulD3Y4v4VCCJni1/4GWy/EQVl2VoP20EKmxXf2P73jW/59MPpcEQsSuWLs17WzgWWlN
LDERYvEAI8wGRTG5ziVsQQmzbDtD+vHv6iFAbSJxzOxjORJCXIe/WDI9W+n4jHQMW1+BNtOx5V7s
PXHiNGuTiX6dpjPWRUO8sf5F2G1kw5hLgQ2MCCwnG+CjeqI4z+36p6A7lOkC2gwEbnwNn8eC+Ml9
9+VrbnZ6DexZgxlEp6RiDqBErx57RJCdWI9NT0VQ3z6loBSSnKSsclbyajfWraJ0mK2s+Go3/bKg
gumxXUqXcAUAWlVA8mzNbYGxkU9bWI5BBAX5yXEqNf41Yj5fQtlS0SBzKGeKcibtCP6r0+MMR2Xu
K86heR1H/X53fLChVeWHTnBFjT2v3nXAhy+6srAc3LQDrUv0VXKqxpWNrCDlDFieHqI/hGY1xVL3
J+W3F/HJx9Fv1g2dMxb4h7kzj2r4rACZVNl1uWLA8rs6lY0TPUGr4xZr7aKzdhJWksTkxyTb2KRN
cI8+kcRR1r79yLgrCUjfFpJ/1jA0I1FMp3mXpb2MgVU8y7lXhMr4POuLMWq4vGX57B8NT1WqNdWj
RbMWR5+bIWTtfjCRj8g1Cww0wEcMAoObWSTQul3dyt4jvMrvmsTnu8iEhYvr/OH8R1KCPqAlJRJK
meGcDHIqDV85pN9XD+pJBu02S6bIh7RJamrSJ8nMs1nsRDLoKhUMY2vVJe+/+1RqTlKCin42GstJ
jkenMJC9uTGOKlUmHkBCuQP/RHi4sHY+uglUO9061zZccopNPz3fNnmMOiG0kNux0ulC1bbQTJeo
2OenUJrhOjwqZjfXEQmmm22D5PSCgwJY7O5nluVHdpON7E6sp+S23yVWG+Go4j/efjprmJJ45gKt
+bz4HHcTf40X7oiMdNqkWRPjC85uBMPfXC6gV/wGGuQwFzM9Ddn01y6P9jbQWwItuArHx56+ErDD
BQ4SJ4S7nVtb8kj7yCSkwyCr3W3YB5jDsWIguS7ayxHGNnsNLazjCeVWY56kZTwzQtJWpSDNKmfb
N2Qc/EYVaGIKN+oRwFff9y3avDdOUfvgIP26P2tG6jgt4kXE7vC43TQKmEL4bR4qkQp7+Nef9x6D
46Wc2mgKThmdapUxHuFFRjaYae07IIHtX+s9KWSaIuXlvFvTFdHCX5mU6HUYa2eyQuLGQwuiwWzo
nGEdECoCgwbFHnYK+DIE+anv/YDuma98BPbgulVyjvwP2gimvYvhpdKRJFcF6a6mWAy187foH3XA
gL2rwHu1zRRMJoYwizUXlQjSuaS9zaHRA2kj7tykrhwc7mw1UPVzsX5FAJ0hN+xnAOb4o2/mJN2S
hnaPsdUpCXz7HfkY5OdyoTIOloeVhAbZZesd2roykd75iacWzvjauSThpV+JKzcp4MzaPOjjAXnS
tyXzGL8DXWxtvAK513Vi9DhcDCmGtFybKnvlre4YfTaI3PM0NvHSrWxaW30icrKCx8Z4KLmLHfM9
RTWZCeSLfzt/JUZNxWn9FsWiHQg1AL/cU/FUFSDNR/iEhp1gFvStC1ZkhJPMyp3WrkNQMVpSnHD9
8ohB+jAFJRtXw+hXn6cAqBRfQR6TrZC7k/0TR9LJeaCPWxHyU8Rf3O09JCFLOy1E+/pafU7PcryS
OjqpUZu9V5EaWE1vhyFANKARY5bn7eEbW3pvX3UpOuDlo9p4i10ppybMqwAP4Y4iZGKBI0xxjGyL
P7jeN1vmjfR+RKA6YbKqqsfNfyPMsNiioVSWVsrRT1ccvaoh6c/RV2dI+HiONPld0PTeb/dNoDlD
5Sls41G0MzNC0X/BuTGRA+p6UYaa7e144lGQCaegBkAFGQrm5rKC1D8EgBDPM2XDWP7kYbnZ7j72
o0tyR29B1e6oHiKr2LOoPh8vAlq/AJnPEcLWfkbI0lK6Y2Y1yL1WpMFwJ8MZ1B/mztq7uGP824tv
i6JSurVMt6+QsVRCkwPP8Mo0m9tUn0iUQ6Yi/HdauS70mi6xyIPP0Ui9LQ23gpoi/P2dpHNJH/lX
eBHkIPAUJkdCJbRK1pi6pHye3c/CN1+pm8oHDYNw6vVHv+8Cs836VnaLXjAN95ZzAJNmHSRKH1Bj
dYY2ZdNkLaW7Sxv/gyEeHpqYPc4wz7/Qbf5TAXVSeGw7CcUJapEjQAvN8pemQTq9ovAtSfEySPIE
F2zAna4XWLkZ0FrWC4bx8Xv14iiYjT7gF1XxIcZzEvWzYP3aashh8O+Ef9p1zWRnj0aC8ZcMEZ80
qWVw6pr2+e4fIIppZGuWx4A8IYZhxJ62z0lgtj8ker0ZizE51RCux6IPLdSGacslyfSUsUEOz7Lz
gbZYjDlux4mP/wayIchS3p23IBitLHdknxPcVdFBj5fCkTssHgMEZbS+nt0yA9JIcbOUs3wPkyGu
WGHsnlrgVIrSA6cwG9gUkgpnqqNiRiwUKfShFMpJO7DpiWexIG7fuCmyLJ1EyEByvUdFSMWSNGOn
ERGa4N93sejHaD+c7C1SQlrtKdsrNJe8hwSALJdDtpLrI+KoauntqANE/PTVhmmyo/NQFHOSoMO6
a2tvygJX6BP9J4CEwEID7AhzQsKM/uR5HBCJXuxCRV+OADRXuPJlTRG1rowBOdoCGrCGy+UW2mKy
OM+r8o2hNbrsJ/L9af0QaKYfkpwMjMospLh7HoxYUgYF/PaACs7UwRpRuO7QVenDlvIHFic72PQa
wH9tOfGLa+EqUgmA8k7sZRv9srLy3AA2km5H3R/Baz3/PN4k+JciT8OOh9INcNbOiC/mj7+zOTze
RnrWwXOWPs9dh00Dk231tNsNVIDPI5W42gnaW7IthAmk0jzggkHMqgSMT0Hz4rL78P1+TqTsl8i7
tLtyzXxTsr2mCSolUOYN1SBt0txsAIiVmrbwVAZmAuqHfpLT9RHMW3WrsDeJaWIY0PfnZNRTFM2t
fBsW9S9msSsk9WxQyK/TdWt3vfyI0JcVdZILHGMG0deoCmAm5V5BdObuicTUxeduRnWIx3YgE1DO
GXF6C7G9kcbZ0DMlkU/AyfcSJTxxr3JDYA8nn7KWNgdb+HBafa0d+ac3B8hwweTyp9hQlm4Vd9Dt
LVJL/60Potph/J8MCicHF0HZ78pF/4C1XRo2Hr5AV653DUUeqaeyueKUncVdko9NxmvIeneae2ox
IUtTyriCUkxfd2yiod6Aky5ppeShnowjHV82a7EMKM7EwA/WdRqIl+mzTo47aXLmNW7gobEXEuGy
9SOg5w1KriL8640al7bZfPHgGuQ4zZTOBNfNAwKLJtFGPzNlfHDw7GjEZCQMYj9DIHfRjhn+GePP
hs1OFFsoirF/TM5yKE9NE01pFAHjP3JEA0q0XNlVnb0g8NS37NwUKPVyLWukQFhp9whs20h82GF3
6x4yc4dzXVeKsxPe4a2zwj8gcR2EO79LXvQg4GBrPaWKMr9pYuf+Qn0ErLDZxvllNnHLuGqzm5DL
fchVB2TNI23L1MUcFos/bJ1vvC37oV+4gR9iOtXEgnqsFYDxr3UwDV4Y6ocjUrMvr/4Vewc4UEUE
ldPvJ8LZXYZc/8aSjo6uZXG0IWF7JBIGcuOBP0ZTplmwSgpyIOs30LlC9HEGP6h17a09o5vhmVta
duuMGyclBwdpDS5BI2MD75QyyqxjpEi4C3UwtBYrmSaoCVyapMqqt0Tjd7u/fMBfttYRFsd51I6w
VgFSGddFENBQkGJussC1X/YDQIhFGM8RQwBdg26jQWnHWZgNBTWp/jptt5kpa5EYIm//Nuw89qGk
3JgiasbC0nkMGsBH5iexJ4rBaZKE5mrFPRljyHTZiZ8GkQpsVYozzB+LxNAeChdON5u8NRyOFGlc
vtJUlMedJ0EEfh/oU20LkMtZvtiJK88TLnet8GuaIqBwbs7wdCOWlex0jUCoJ96E5TR5zvAn2Vqz
cJDf//iPPOkp7ZdxgewSJuKx4pQkyp5FT6VFhmE4/x1RQ0Wflk4duToc005BspTSIU6705JCz6tq
i8qPNc33dxlS89pUqNfvIs8l7crDe34iLW1IZ9N1E0dbS4s0xu44BScXWIIiAvqdLsuhBGWlaOZK
IlSJNdT+j+aENAcvRnCagYTSsWUoLHyc1ed5FeA/GGEp1+mW9Tq8Lt680qQANiZhkQPg0i43l8fu
p4TWBXJhlWvFV7Dyzj0FFfX6Wf7dtDYT4U5MpLWFSDCE5bEYDnmHrw0uquaee3+zCqUMoMbHI5DZ
fGhOEkc4ajaSyOUdHL+glLXJBZfXI+lHoB87AmxZD/5VOms9bT8wkSKeJJyJAza6xpyDnAgusxLj
1iO316HPYFsupAdfBuwblN7u3S3VksqwYhi3uXkXwzzP1cnr8lEmcgq7Dn/PvXEV1N7xceFv/W09
aKadmJ1KD/PM7ags6KZuuRdvsUXd+WK8kHVEkZQUAJgP7gv3xkAIco9F3AvElNuToZgS8MH6HqTk
ZaAnGzNQP3L8vmM5h1iWMx3Hb5FqUALN1LMguSiNkSgs2QaEmgpK6X8YP4E9D1ZCrozeISHY9oyy
xgCXca66TieZNZFwUBhJPNwluPFuw1TFedpSyp5HkWqZq3IPixHI0bLB+kpk3PWtT0eRNBGPz17Z
H38DLGdISQrb3TL4MrBs0sOoFR9mmmJiXCTRXXQ0u97PZ5II3inGxmT9unF7QXTF4L03cMqKNG1P
YM0Kz590k6212d85c2kOdUlVri/HqaV9XUZVG5YPjsZntHyg38nJbbbtajZGNUa8kvuUvYp37xeq
DtXl0DzotHAlFc8YtTlrHIC+iorj8a1OA4y+fDULVZ4l/23JXc5z7wp4sf1GcqIZmN568KNVusBm
PsQBAH+nvcha729bkmGHBLyWY67SUTXVKQfEbGGExN2mhJRtJVOT+TcpIYMh8BLNGASM9TsZNmD6
toaFMS7+XFW4aUim/hBRoQNjTGD719TwxPidj4OC3bHNpGSzPd+UQpG88BwxhFdfuNrh0zJTmb9x
1/lBytf0PX6lFTzuQVKkzE+IEuORYBEZVf5BoleSK6O37rI+2S1zxrASy3VYWtQqM6tKdV4f2eCp
yoRh3ACqptPjupaRVgBLfmcx/dDN7Hw/FbLfkl9KaNkfLIQYm+Xl1sVErt1Hyk0wWE+yl4EoDVIx
bucWKgCTVoP9CXFFM0so/zWmLKR/9oi+ZeulP4OmmeJ/JBPh3JdsrwqgT8kEDCZYM/FybU3GoIkG
zVt3N4b0jY1nXv04LOQf+Y7tAkyDoMgHxB4DuPXE2QiS782qfkFZMdpBusudTAV+iYFInt6oeUau
bYl+H2N2k5v39VaPTYnNgStqt/+dxOZ3dYnF0SA1AEz9aQcaf0qgSTJ70BIeQas1i9ZiDMSVfpAQ
zj4mZ+gscNIF7m7cO3fvApfK/nY6N/8FYTHsNvgUANJLdWJ8LZ19SU0mtkFFy/0m65v2Dz24lHH+
JVOq66myfk3YpsQJOKRCniA9viKZku1SH4ot0zkDt+xtwmluQ1WQOcDVjU2xO6qeWNfq46t6oxqK
wt87Kgm3rX+l3iaS3TYd1rqRGF6n/3/wX2JnAdNLdeg2YJauQcSmzwmxTuP5ZkzqEjqudR87T7if
YKcG2KHJ1FRwECE0D1Wm2yFJYB+kDk8l2f+xTNSQ6YxWYPAuyOW2aAjvrJqbrdV153GRrMztnxx1
8MJuvf66fejLx7xUM9y+3C+1+0n7gIjVc8KQFtuj1YRmgqtNM8rI6lGPX5+mZ3NM4b6X60X5cKLN
hfySklbEsd8GLFuUbVFhxOo/wG1pZjb4VxYeQzi6Owcp2w7rjOCLegBby/iCG4FoxQh0AMO3bUU1
F/lMD7ARe495RpywKIepxujEDwGGrjBZcfHl3nL6BqvWbwgHludaIvXhZDEP4K9gv4CxbEn36EeP
GSu4xVKRMoV6c/hohMK3dElmy1ET2s/R4zd6V38clFWmVQDo7LsR8CIqIU3tEg+nI3tS0T3Ih+Dd
cCu4Ig15j++hJ0+kP5y8evuOSVqiBaa5IfhCWqxvcvFSLBK/dTcLhhjuLAaR8o10G3G/LGcfaeTD
SHpq1S3sS4x87YTVessGDC9htKliJ2z4zZSUuIzHRBVZ7OOHuogY2u55fW4kTpoKYg5M5WrpE41/
5tg0NeO1tQeMB1XIYbu6GLTL+QL6oQ8PMg1/qFn0Puaot6yE4VQ7p6yhrKQH8Iyh15ENNNZYxc0r
JVshsG3BLDxSxi6DUbsYZTptj3k+bcUuAGqBBHKCQBaF8f4logJOBTUVO6QVVXgEFyF3FpphtIEW
y0/B16qK85sZNHE6K95NhvQgvjFab3DgBPtAKDDMrnSKp4KPkmdSqHyMFMvp6tbL0wY16iEwLy9B
TEKqgO0GckQnyyCV3cFtIc/OtXmtL/mzqZ5+Ej1zwDCWgOsrJVWd6paWZ4sQ3y2R4tcNyX3H3N3K
17NkQ2zjiIkS/N7Zki9nZpbnYKB8D5ihVdXp62IDczPPXo/fsY6jbvTbHI49K88trdr0WFh8sGX7
lVHVisbk3PVgl44bV180EpLDR5bK7ex/AKoZw8t+G/EGlaMZ9gyq/GOQx8n/5hFyzZmmEgnxU1as
u44wAtqgHxmXcHElnjrH8S5p50hrXWFow92Hfx8Q3L3mor8QOkRil79GUfr+GH/N5VZjEO/A/Lhi
bYXM++Oqk9uJn+a0mIVz1BIT4ivBlOPK+N7rgLbAxS+xh2hkLbYt64iG3nuTfQuITzpuxD2x01BG
qRxkGTzrTeoEUH4FJM/LEhGuQr8b2SnXaCHJuqw29VP9a/CViN6Mx69eUtKRZg77KSKVO6XVF+Ef
g7GPGs2ndZXU7pq/yf6yCsUF48bma/MkgiwlwiZTNq6xf0r4JtJoePnTgD6NZoZCuqXqxf3KBsPv
e7lyhid1m7XaBzzi02WXKPs2PNKDsc2kAP9OWJrGCMeyQpaPtECsUTw46Iyr9yuTENKYRQiC8Do1
FVDnHLS0pF1sJj0KHoWaJSRUVh88vUZkHN7VzxQPwlTR/gbjW5dTF2+dudSmK+ed0+IJdcCK7Ass
TcBIateZUvSZ3eaOiDjGsnIes/qj3n+eiGDzI5mjeer72+5EfmSKC87s9/BcM+8gkgCxLH4lDZTw
h6HWyBlS0DzRRkLArrNjutVfVun5YQ8YZQcDpU+OnjXM/M/Z9GhFXoDdPJW5UAwkca6St3YjUf67
yAJ32JbJJUSLSlQD3S1UH0UnXcK4cOPkYxKnfS/jXo3f5LROSUPvI2IasIWAVL0W8lQDIwOk1yW9
FB7VLr5+8DGUpqpa2zLhcjWpCVem5+3bP3gT4J630n+sq0uKEtX4spzrQAeo/CPnfMs4XdW8DpCC
IxbbpAJziEiEpjwIph7RO1H6IU+MRTEiWoWvmKLhNHe69C/UnpsjVFCu0YRoW1U3vAPMHDjJEzYH
27f06wgJA15NYGdsWQPS7TGYpScmI7HVh1Vta8Y1jLIqtsxnZzUuRGwdTBpRz/KgO4cbJvjTGMg4
Rbmo1M5Yit5hDRdRZCd9Mr0kGk2dWzR4KI0htNdpN3jrUgDS2is008R5f67iWdtFbW+20letXNV2
emEcuFUxA+uNP8GchnaTZC4IIQdNUJlImsGbTXphicy8t+ac6opeLL50dRrxRszijcHcZf1uPiPu
5zC/eY3gMzFmeUQBTDe6/wJdyGQBUylXuzXjetIHLI8YdTJxDq3hkdSgt8YWEeRSNzsY1/GLpIJk
bTuptt8HDWDskH4ZxYHp55S75FeTA91poX4MpVteCoclwLxuupIlD2lRrTWod6VC3NuJvnTqGk9o
OO8Fw1XDiivpPCz8Cw88N5KAP6jJByOKUkDTNyT6Z6XyejIhTJhnUJI1jn3tuNqTHLSITRZ7ush1
BhzBE3esynCnJkUZ7ZiTljldjyfx4BGIv2hNjdrO4Bh3ro3+HeLx0j2BUifwUmrkRpDeM/qP30DR
xCz4ttLI19d8ioEU6G2h30IgtITdc3BYMQ3jSdl5DTVZRgAZ0oefrgbvJVA/zfwoiLNc7twyrZEH
A8MJlf8T02zSEjwyguq4kHfHqhwRaf3h1KllVvdwPRjGLyFeUGN0GKwr6a9t4vdDJuh+PiPDpX6p
AEgJt4mr5mN5K91+yDH1qV5VTqEvHuPlvO5qEjaTXx6HWi+JVadielq3jwwQ+4B/ElR2mCT2b9fa
y80URd8Yx+V4ohdkuhJNSWY9TByz71x58gAQGtk3XD1ujjjZHfClUU8+fb4Ux5CvHLYWeg7Q2Pf+
J7RLG3CkYwhX04w5tNKxpSQif+A48n0uutQ9MBhoFuOzMzfRpuhxgzBWUzCUW6YErJsI44Qt8FyE
gaSDoI94ekG6VN3P9NBMTM08yk76FF3H/Z35IsmxqiyhVUN/CXc4Q+tCP2quBynNt/eSFFOkg9bG
zJY9TXwEAnWU9Q/YN7iRSZLHClRU305Ikp17TDj4A+D4Ibs8Y26uavGnmEHV5Tm7XdDk2O4qpwvw
fbP/FnUaD0a6GVNA8TKZx9O0Lm4jJT30cOUUJ1SpIgCdR8gFvCPRh5V8SwfaKDcSohJCWnFx5xQl
CKFkor0J+3ZnY/1hxEEkSOZiEF+NxSky61pRMNsu1nv/Y9czh2/tsNgQdQh9dNy/SZpuPTh+a7MB
p43g28KsjNFVzqFjGwcS+N5DpxF3cF9+soS4uv7MUXnadiMj8SyRZoeyvWA5liveDpcHg+wH5AF1
KC0UyxnUBIosGigei2mwDG6ktiA+omGWGlinqrfrpf+g0yRYNr4OPXxyk5OpO3x3VnqQJ3LjujpZ
2kjIIn/FKnyafiPBBfVJAVgjTvjnDEG5dnslAsajeHa0Jyzf498Ylc55gONw1WJepwkrUeU9uRZe
RE1QEZLcvd/XNAyT6B2EQaStKzp+tWZC1PVKZfmDu6UjDyOBPcgeSAzspjM5K6dNEJ+oRuCMTSII
B+Z+/Qd+hLm+Flfn5xvLyhhsZRgSCHdBPhDT4qGMpVbYx2/8ck5MaQF/sn5nwxV0J/+d9YHQPh7n
v7DjAkv711DRbI8+N9EMEl0WdV7MzlTJwabTQGmudLnsDUdahnfKStDMsfT3aIZ83c3nmYSX7Fp1
+a0JbfAJyDM3wVmB8yM0K1FxrV/DFq/CiPaO9vLYnaO43jQ6YBxS6zjUc8aMXhDOJeb+9gmUzhcj
obi0ToQ8hPvVgPkfr68dB+93KQyxrnqt4KhH8LigDUIoocnevf8AzX5haV0dgVWtU663rdobhLHI
/8AepLWWnVNphIdoyU5XsNXcGw1ui1yUyT2Fj5owz9E3OpM7HgqP/bqCQjyjjk3xBvrcvlwIzcAW
doJaRE9uCwOP1liR0zKbHfvk0bRckvsV6ioHmetVGiPmtuiMPvGBHxXmzlLU3TH/s1cBqZxrP/zo
LaPAjVsf8CTG75JoRxUfCR8y9mCJ6Wh3OFPX5lptd4po+9w/vboea9gnyKJzmdKz4TF7kJwE3U5S
yl1FDJy0jXXUJwEcI35I+vVq30aItMyuxt1xwNADToVnJ9hFMHJ5206EsM+1nEz4Bo4ctK7cXSY4
KnI4waQrKuK/MtHizwSrFWfK8lWGhYJ8qsqW87zKPt/OcdrHZlHG3QdtYnK5IvHf8PMmUMEgIzGP
8h/JSEaxP3g7tMHjBQ27Qz9P3iEZZQHMvpmn9vKQlAR2h/J24MVTx31txC5+zsmk8njb9S2DYwH1
KaPCZvYjEPhATveHOc5T7pjwICWbwY18yxNk/HJTXb1kVey+HUQBfQCTrBfAtGETy7FjXRmATB4V
RUZgdPf4Ddmfsu0Ed4rqSlzGXTn8v6DaJCctPqZKmbaOi7UAh1SeBjQpqmML8hvsqunOlCoTBAH9
24h31Lsp0f6WFxZOKOUkHwjbxO71Jd1tZqgHtLaqMCxRfhRztzb41Co7luSLFVIb8/9ljph8x2IJ
VrZYl2b6xJiL/2/oNkbS1+5QeecK9OTDsTxNIUBGKTi3F+AxbuxaTTPPqfePDiAemtYOdOv5pzfI
UczU4NSKYs0jaTYwB4x8Z7nsiebNSUldId5vLU6c6rES9bXK+ma5x+/6EYY94BaHB95FW6mhycAt
Lhr3IdjOMbUIV0a3A3aawhvjWGV1v7QRvqOj0zD+NdFWH3Hd3Sg3KLGs5NCllC2CqsPNCu4J3A/x
lt3mYL4c2CMrFCvtWFN+9pKbTpffHpmZ28nXT44cy+8nH7HTZnC/5CFvWpFBxxCtjjaA93ev8QuP
Vm29lXZ3FBkQlF1Wpr09sh7VlQHvzA8dW/5n6ydEFfom42k7iudy4pwMsCUoo3wbQE8wZ2/Lw1lX
fbjIUaGCTI+c65C/2YbUfIf5s4GWDnzrCziJUMBmV0tK1oYViTQ/vovgCB3Eyt7BKH3ubM8JfScX
f/qCHDrWgZtVMTj+zy+HOSGz3udecNb0CFHHwP000LJsDsMORmMHQcWQEo1Y9CKGRa4ODJeJZCLB
MwtAQc9uq/q//2caYN680vgu04fbzxz8yluMTAY7zP15Q6+kSrAMyugiyb6+/dSId5fqsc2QRJl1
5XEj1mtjAzMpXxoXN3Fs/vBj+EVunSw0u0PuCThz55Cw9qc7l2Q+4B+nUdTt/B9VA1HspTfiPJmd
nhRVP2oQ9oZUIpS4dTwPFQO0VnlCmaYWWxmpSvhGBrzCVSzJTsW1bwaKwHCKNNBwUp0yM7xmhAUQ
WWKuazZ/BwZwTJUYaSoDxeTdzab6OwpwRFFXazgmZRni1H6mi5CLyV+XAlijxaQe9LEvC+/hP2fJ
VxUffH2fEJzcgu0FoqCqy4Y2eE5U/x8zff/CZwrxdxme+G1YUQ8MNxM+d8IzN5JRs5gV7vFSDVZ7
dQ33yS270CwN1ngX71Ov+UCFD86gxAol9Ojuw2fZsJ25M4TmIArY1a2CoUrEYkXDemvzarK1yF7j
7Mhoh4DVsG3du+G8VJNWWnbWhgK0y5S0pF0g8je4OX+WLiWW0JMohVrBx8V4aAXbeZeCRa2K81qp
q3LHHj4XftgsNsI1H7hI5+PNMrEEhEGgQquQ0OGRjNz4mjomNg3QgKF9yZoecyOn+eR/QfgRvPo5
EOz/hH1EyH3GZtoZmW61LsweTUna2ehRkEy840zJF44/vRka4UhijVrWDSTGkx5Sj5UwwVGjH5qk
vP70IU2oknZPdKF59m+jbQr3ib4B1vqU4SickZColFoCnr/bBFm4cA46NeTRT/0Hdq2ozrn4OzIz
Lh5+ktSJuRnMjqRvFbiUGFylXLIZsytB5BuM11wcdp2LMtpaVl3lLAUwDkrVFlckzF4vD4X4pHbs
ZP0dFXVQSiZs3SoSiNaLJO26wVq2hff3Pa9m7Fa9svfh17Hqr59hNVvsDRQIau95+RBSXnLXBxl0
/+xN52MekbohzrdFzs76lrCHWwMJFoZ7/wLjO00IgaQ4u25D2YbfyBFyD/tEonEqhid9RrP36qMM
IoAlmG89BUWBx0S8YqWwirlSLAFECxqS4zmNG3K4DaGi/HCwYmvDHmAHUMR6TPAl3oUwuwXM4gUK
cFO+8502mwu7n03SccCceVw0cyPYQ9+uwpyMSmjZb5bXw3RnUaVvVa++VqqWZPNNyfGMpVF2VyrA
7Zf+wa/Bg+uBQC/GLnVhx5AAcmh4QR01qprh3MKRJPSn+5+g/nirwQDhUQ/WumjYa7G7mKM84Mnp
yuZd+2cqd+V7AbpdEBhH2GlHaXqh4SAS2AgNSjRF1w9N3OFhOeKwN4rsswlIGKRMbpNW9n9+1ycq
pi/IECA+tdovmfQrVaFSaKiITLpl1lGRh5mAvmnwLpmYYMxp8ZOalGGZ0jM2NEouTcigI5oBDKan
DYSwDUVSDcLdKK9sM802hcpqshJ3gz8v2KaCc3QXEas3jc/R1Ib9dqUyHNpMwgKjr5ykktnFq7I9
fGZ9Pp7+RTz5YVswTvzOurO7FIM7IDhfC36xcLB4d2xE93hPHntaBVIjmXGXWgxNj/HS7HPgxo3j
JReA0xEpcNIyVAW3NaCWS4rtDkeWPU4P3NHCedXEFhM3hc9s0HC+8TU8qSNdnEhvydOwJKB12jiL
g82LoLtBZA+XXmp1ogNdu8RiKPIn86dXvb4+YsZHyYEf3Id/SDpjlQ7EuOXhKibTU9O5MEj8rdo9
d9iWVasN1rXXj++kwNh2FMqhvCg3ElZoqbLdTfskRMBafVI6uOMMcgSS4auz+LNh0tX65+8gDlaI
mr/WIRROu0G+CLFygBL+pgK4ExhnZ1KF2C6DQFpaR9qJrFhIMgMo+4kLsPX+INiy/HMu5IhakQQQ
mR4qvDqd9WLtOAASDZq/GcVpXaOt2LYMWf14ca31TbKm3POrsw1oCD5FNJr/YlMhcpq/0nDWcWpq
d8j5Crik1p2NJ+JtbFbi1akIxkBzh+i3+41WWaryIydZCfsZZxBin+SX2n1bou34W5yBsic1qoxX
7HMBCND5ppUtqK5F5Sl6Lfcpyu8Y90Y9mGj36X+Xcvxrv9IISR6LtRGcEKIYJLmdBwtoUdS+SM7S
t0eckgFP6ND8VwtsjwlZ8sTrkLvPuXW/DATDrQAl0Ztv6OB7FArz4aAA/LpPatOdp5cEUAdG9Qz4
VY75eyDc8rHVyJQl17nFi6NtW2KIliawptpmFRqCsy3tKPoFs7a5NXNxGiA3x/G7IlGQ8JqwsToI
9/DBLKt3ViEmoXBBsQP+diCdHT2rhqPsNz4JjzmsGqd5lFHdhEPvdtkwhViFbPCee9NYwoHoBVK8
kC92QIfkPynPE1DuVsRHiISn4K0Jv64oJofZJyCE/c9fPaTVQ8tzEMh/W7NJYzvTAfbbCwcdA6zV
y0F3iZjY6M7CT2HiFHQ74OY/ywnQrF6ZyZhMtT42lEYEdkDBd/9FS/l5PpifoDzjd7VuQncurRla
cQElJ101p02PB+lOyX8mJGLqNlkZtvOx3mRM/mmryenl3P9LLVuGbFZq43c48LxRo1ysE5cW2VOg
YGvOZ0cf7jmE2eq8pMzLCH8+pCBg5xyaJmPcUfh6Aj6jqal6N/AooX6d3H0mW/2lYAjudd26rJqB
a8N/0Xt/0Di3GJI4ODYvxuVU/wDzCj7iSg9vEeCWoeUXfqSV1F+/ejuCwJWHC61wrccVuJ6Gwrzu
AE67mechbVadSQutsNK2vxw/6CrJ4ZD4LNR95z9AAAEreChfw00+AiS5k3nZx4XCkUqbiV1ZdOsJ
YFnjR4iJwtS0e032xJJ2NVnWbcAwNfZf/ol/9Zj0UX/4vz20dwyxfbL3xAQkqm891DZwQ7SmK8e5
DKxBJ0uiE9Q39CdIAArfcNXs+nS470xzHqyTaD6x33Io8H3736Ku30gGzJtbKfFwI2PLFzK3AE9j
aA6ScOaru5quYIBSqS6/TpUqoV60ZuBMupTgQ2X/95NRdCU/l74BYeEtCbBXTKQeSTnwtp/4CqZK
1x0ebv9OjnCx57giX91vp2kR9Qmh6JKa8zEmyxnZhb+qSJ+QBmzyTwr5uzEmgjFnbCFX+Si0k3sS
zqyNrBdcbWj8WTXZewmj8UvwrrwSIIPCT6/CaK1xbfOE2qfiuJFijKHLBdzJdE4jtmYlegS1v1Q3
mqWv8fFy1XWhM4D1zWnbkzMG9bumeebPzerZxdjAi3f0ot/07UwL7Fh0S/ciMlvtc+30O3cKgMy6
B+fvhkpODSS3aL8/LPUvy3SujUHYWDQnjKnlVIOKKQz1NSjM+RKfjXjG/kaDTtosjX2+2XM8IOxG
NPZG71sDh39uGkBYP4P0FT6HjyxvqZslftaoLt/vv2d3T9/82la2j+n+0JimMe8F9tvge9WakRWP
Jr6A261fuAo07HaH4b/3xQI2AB7N4N4LjoMWjG8B8qHLYH7gGAZocHekWRi72tudYc8dGjZNBs8P
mvOqJgBIHIrRe2OnOYOTX1ZG68jP9OlldXo2X91k/faSLCq59AC5es581Z5tzVTbJvP7Yg3RS92A
Ahc4RZUvuuOwOzP/DNnpthsyNAW6upcOUMszJI88pEFZWeo3MDcjWngHXYkNBOIGmBi+odyscYaT
KgphrNud3ZAAMnFDwhNXe/q87++BhSH1BDGL3aOrXrRGmbRDUwO8cwxOpF/krjP/qcJCLUOGPB3j
2/0ivRoQ+EQGI8p+VEvpq/GpR8D121l4S4evBAHXuBus6CZaLyy+tg/WVjfitCSlPPH+qUnatk3g
CIIqNx7fbxCWqmngvJtMZHdf1OJtL7ZVNFesdiUf4/CMEIp2hQ19CJmklrziwtR4hi5B8QqLxCEx
sKYqbL4xaKktaeDJys6cMUjUDWfbBYfdlD2+ax8LHzUSbtD0AvKaUKlDjULI74sfm1Eckqh4tkAf
+GyBzHslzDr6pfw5BrRHBATP76Vggdl7tNjfCXzZXfkOeC1uXYA2gWa79eJBzskxCdlgOirxqf+U
vbtc0peM9wo53NVmYbiMKHpBnlo3lYAPjPcIsC79lvlzKWyf+GQMhoNsyp1MXHTGGSJNUXVHaOy5
WzM90HPNzz0WpD3tN0y+2qVI4tZN2PYhO5XuAA5hGY8n5vjgqk7z+Ej4RAMetdrbao/6ySyHyjkI
UH6kgo3iGTdRON0hmaLfAnaDWkTFVLKT7of9I6YjW5w1TiUKooGtoMjKvfJLKgi8544Y8M1l9z/1
KyVhf6qdOUsJx9OUhjOlItsNCnmbKNgcG3abkAFF7qEtplJNs2Ye3YsXKRsEUQbKeaQxBrfchxxT
VraIrigNUMaO2Esk58DRqL1vTXPUNqYz9/XbMw47dLhIiP2xaC2suHSrzZ8WlUKeCfrTHtGtbkaM
wzaHVmqj5mBgZzfBSxwLQu14injF9S/iSH+wx3VyKQ3Cv5cyYX6VOYjcLAwnilbFLSO/quqh6T1z
3J/pDsLtOr9Vc9frOR6MdmApF/DZlyu3tjd0GROqXndhXS4DrGQ8LFMi4vtRAcak4B7GStyyR6kQ
h5x8oQvPk8+k60Koseob0acNYYbxbqPOMhfezsTvv8mtLtCF5RfcWlB8feahorXDWi0Nuh336oMk
xjG8CHlYrPlycCqOUo65COA6zPcb+dijUOkOyBKL7ziaR6l1dfE0Mw9aHUzwRFrT30JkeGBRejdO
8aHxYwmW/L87VkvwL8M2fjQFM3PDpQuzQNUxkyxMmOUnMU5LCKA4fRajsHlZuvt8WbbKYoe4bTxZ
k+80KAAh2H0cMjMWlHJwlrhUUf+Vt7W3WafQBMZP5tIuTDZOrW9uuOnI9iYEkpu/Ha6Hu/FWgXjk
b2juQ7GOlyLaapUfNqG6OoBTvCpDl9Xl7odA2H+dHWutqiyM2R4TLAUpREZi+BvTy9IPfYCP3xBE
grJ5/1FWIhXNiLzrvwoz3E0TCA+ZfP01iQ7VtaAMWWmnzW4gWhKFVnrTZfp3NSi9z6g8ZBiPnhlw
7CViVg62NRodguHMC6R2Hpd+WRhsQeVnK0Z/KKd3JZoyvwerrv8OI/tgRvjgyGqtfeR/evc2w4+K
/EdhjLHLm1Rva0zrueMY0NAzgs/USAFjBjFPqEBWN+sGv2nnjp2vAukx2uQ5m8zaLBzjD6biztuV
bMSe/wBjpJxocEE0401IjH5eGLJb/RSi98St2kMT6sKoaGJR6T241TZv3xI/PjLp8o5IHKhM5cOh
GAuc28xodbVsFYo9rnTjzeLGI9o0QCegRDBEJbKoaazx76o/QhqheTSMZv9DYgeIf5xffZvVLZlg
Eor6KYzMVSPToXu+1uW5pDNyZl02noERca2xGVhba0IolGkfWW83jHyzgZS7wXlNWdeEDi0MM6jL
AGYLhB6rFdtVUcYMo1/DYLsq+XQInNIz/vKNTE7SR0Ozv222Gt9UAsYlT7WAmO2ODAZ8Ki65PRQW
6RS3PaP1qD2NckbUQAjpwiueZGgmp+hdOlD2NgNHGg7kBrv+ntMHzPoPj7SeX/Ul0kK4brUcc+sF
Zmbtqma0yDkGlm5nhqYRVSDh94x+VS9Juhm9SxT05Yoedm1wU1t1P+lwM+Pg1HoEilr9dH9DrUI8
bI0I8M+E3UEioNSwNUqNkNkZwRiumGl4daNbIyB4XYCFZ/yyDH1q6Z1j/URNG1CJkh8jfIvJtz0p
XLPmXmaPhF39FSQ59VXVPIx8O9dTJ6SgU2UtmQYM2c2ixDI9GjdUPPSLLTtpf0erNmBIfVt2hquj
CsnqFSYUbQFKYBYNmAMmK3NLQkE31N0SIUWPih2pp3b6T/YNjP0Jj/WfcyidsxQGQFw7Ax2YErem
5L2SiviQygNq/uZnRA4BL8JWgKYPkM8jezc3Ma9XzowN1O1EIxbzrPmrQRlc7lMjs6+YvVI6VGc0
q62Qq/qQUAYBOyy+MFanHPopBazKHNniyp3N779tGz3460hw88NfICEfiCigKKxQ7FtSEXfHi6+/
TL57Q4B615NKILJYThepT0rdiQnbmnLRt38slXjc3zc/H2WG29ooeeJbXAWNaszEOEsUxH3IIt8k
/IdFHRa/hOYKfkrPsoIkkLm5AO8MVpPbVob0x/ZqQbVI19tP8gGK/ZCX4GGalYFD5Lu1ph5CMejP
HjYxAQKVbRHlMBFi9vwtgC/Gb3l9CCOrbPjaCTCrc8AyXZN3tZaF+12+Ff6Zl47Bi7zGzvYVe0qt
aFzfhk+V9N5/zQgnv3eMsclNDH4GdS6F7Q7jEyq1TVzReW/A4+bLghUz7/PYRTh0VbJCE3rvqZYI
/oTzQt4b+csIir7K8uxKI0Sinfv2HlJQ3NyoQooArKP3IjxeRoTE8Za/y/sPG7pwiAS/GuZ5BlAq
god+jkISEb2nMNH8bRHrFXjW1ugbiPry/0mTImLuni+IhkhwCl7V+r35EnuHLfljVd2iL6nR0BG3
S1FkrNKdn7jEtKs/AuOD4waZjYGwbDouee0p80gDKKPWTKBwNiMZkKKwv6XdXiw2IV9F7qxFjFTP
aysTwmo4Leo8wSx/2XXcr4ymuXpXK783XU29AH9UMuFCP2juZ1p0+D1dSAgrz8hs2B2f6aJr1XFW
6B6lnrh/d9YH//RYd/UmSbJlFRUVYeyqvJ6F6xgHkn+Dd2HDfAvh60/tfRBg2GkTUwH+V06mOcJf
rxruFgTCdiSGErCgCKncifs5P5BLwFKfeb9UPQNHabEEBJXRs+6sP0N6IcJfWB5YEXsBG7MzK0eg
LOpUF7Y3XZgd+ZLC06cQPnkXSfj0Zp+0QKyzKBtAJtDg76DeJv9k/iWV7a7fQYgMOrtsfC6yxOYL
/PvCW9LVzCaxYjVAPL9pxkNqkbC96hLtRgulgRbN+RWzYNwG5gjGQ2XP7dlWWwYGmHzq8OGmIfqT
/k5+iupZdJhIuTx0HUXFlnuutW4Nei5jTLXsT5B218BAb4czVa4DV7ot4olT2uEw+E6wuSgefblV
tKXySJCVES9/uhc4XUnI+HYMQZoqfhz3pSR9O1v7payLZtyID9BuPE2ONR49rtEHq1w6IQDTE7SC
UgzXgyL8+4jyaKcCe9Ll8fNZNy3d//EoSggeEt1VAeQ2NfI8QJSWWG6FqhMUIM3uGuKCiyF467J3
s/SJZWaJGqYL6ZxmCxsbtVHRlS1qCasQP+8opD4HlgHIk4L/KWKO/x9554xz713D1kMRDmp4m+6y
FmcmA1qqXo7KXd7uAttPFgdLW+gliT081NLmE60HnYVd+V+64oP/u9brjH7H/qxFC8Wcuk0wScmp
lOxdJbjmINRbt+WSO7KOgSCgIg4eM+XdIKKuhfcy5FOPu+Z3aAbYd9A3zzi6tSI8MkGeM60vMJVx
tnR30K4CCnXeY8YTNuleLfM91GWDhA6GYUeEPRVeiF1lfZV6gB4EU9AozEKAtHqrqkaNCJPmbAFV
JMaXPLkzM1/wWUQ5diGzlotYRrAdS3nBpuaRWxUzarLbHBcpYsGj8nJp1uF+Fe3zEAnaBb08Kpkq
E4mHelfiFNUyBGbj8i0ei0CH9OQbjuyvZtWUqgGaaGx/P6BuxAt/UjfIfVD27WONGzantWBsbVcT
pHwgHL8lCy7s3WPPPRnLe+fFxtpcNOZ//dTc9GsUEri7k+yJIqTeaJybAgZHDlA8vzzMZ+uH+Vep
XSY/7rHnx/ufrRSYJYrlQK6vbGjU3eMVp31Xo3ClRFwEUq5nA2+5de+RvgXYU/TKWvmcA+1aAmn6
ddfIu2kdBXlrdKs4/vfrZPdSzg7Zo5ql5b4Wv85+h8gtJEYhANrwo9qYPIeEn29Ecs+MHyg9YY+M
EWwOaTxyXY2lnTNrrlXJLud0slTw9Q54pvlXxR+k1DquDyeqTjbhONeBXlvH53bjNtlomn4ONI/t
1KoekK23NJvcb/yv/gkDun7Nz60UQydhTfUlowUV2nnYBsntbTxmFt1NsEX7ScIODzzSTqN8QATt
88S6JneqbF7CQaARVsWzm7WaYIhAN4Qhl007aePHICXInPX7BTL3TWhkP4tNrWi199+NyXFhGx/f
GePMDR2kRuNn3hrnwrWkqyKDh77tA+/bSk83NhbDYOWPubUFwWLwbsVtjMEDsMeyMvChWX+ClmrU
aLTAVUiZHWOMUs9sT+agGsshLCHMWYVUWIIZ7KWhhqhMOv6Vw0QfqgpExkDkgRL/uPUmqJL/Oao9
Zwg+IHULbFeIVl7pesEh3I6iGqXlYfg+F9OQLyVc1UOPLg41wp9eWgQdsGmZG0geSMsbPha0IYT0
aYsc7LFfLnTh+YXfHuNBoX199/JnMxlUkF1gMxQ9BS2vIrnxfatDOF+fwV6fHKSk5CgiRbvvInzX
4Uyy1p+EMHjSL145h1YV5wqGVo7lI6A1ROE8AlHnXH6eUDeH8bpy15YS3phOzeHW/M0AeaHVZzl6
wHX9WivMi/8DzKC34ypxRT3l0HcvCNHzBRFTFr3qowAxScgajfjIVqKbDlFiKaH0GpR71P/2/Q5S
DypCNHgCUEfdPsB4USE0tIj97Gg5z3ESzjm0cM53DmlFkNnJDIvzkXYsH6JoJjVFjApZqVy07/2M
Kj6dEppp7HNRlQDZoLvOYeqFdtDFuJrnx0iVxx3munk/CbbOOUx2Hvqw/HrpEE/vmF4kOdZbOB9v
pXkArRfJTckv+meK8aku0zMi1NVMiz4aAvcMBqCb/qp2aq+2jsghDGqzjBjvTe1Kkj3gMOpEY3Xm
82ivU1okwnbYRleSxJgzPoLdkkbk+Ti31kMGvWX7FkXzOhCtGcj/A+Xn2cr9NL5SJFglWc1WuEid
B93C71S3blgFFphl5Cubqu88HbrB0BOjmVHAR02Yg/Hl1MDjemzRUYQcCb6VHgcH3jqVasu2UsXo
WGxOYu7yRNXr9a+j2FbwqIEATfOaFt6jJ4Ri5RBxVfJ/Dk07oZbcY0n042AUufXa+Ak7ldZtRvvE
6+qtOPpEoHvZb71Oq9qykRRzyJ++JCmc74SOgtOJBB0Zxv3C3PBIAxs4bwv0WqT/U/bTi1/Ctjb5
KlmNaOTu2XcFwKBDsKg5p/xu0hhaSbR1RpHms2li06CAf7eS+rvkiTubuJou/Hw6JXZM9Grs2JzH
L7RZiQbNg10OrxSqN5aLxj6FHR0SrlTvWHBQpKa2fM85cb3MTS3nhAYW4ysXfrWxtWMhkMYMvAP5
mpWNyNIm+buoODmJpTmYqJ51uNUD5lqeIunNutYK7501EzENHFG0xoJjICAqVcIgm0BrGU93P/0X
fq6m8562KQznCu2TQyb92/VDJCQZR/AlE4HeP4+uPMdqTAps2ZWUAkKp8mKyLmIuXvOW3/jUGSIx
pFYoKxo44ukVqkSdLOXgxI2hwlDuxw8aRqRccq5gsG3NnSDmPdQ/EytpAqi8CY6ljDd69gSF7By+
/FCbbtjX1MyrqTjHbQClKfrOcT/IoH0xgox9P0UfLw6YgyxmlsgLMvLSzC3me6GzJ6lOUSe/29jk
/hCxodNqdkq3MtF0ZDuqQSP1jN2a3gL2nFY6BmTnlFGMPLQIxPtYHOCU4+Gf3DpBi26BypzBDV1U
9LATreDhA9YvfwyX5wfIMr65dSt4gzYakTHt7RmXOKo20sU/R/7Ns5v6GUe/NqutMjzq/wLsNq1F
I0Rngx2egUH+sUYx+ZbpgvOGNNamxWo07Emh5AsLQwOjOHSxxVUtYZ6n6RcOS+4mEqGqM+ZOxBWO
xZpq0WWKuqXYNllSDlJEFUS7eUkDl6R8gb5fDOlLettJqHv50U/u2LhpuixLvaiQhqzSrjdTg9a3
EYBIlfhfvumFBHd93zjuHAqcXfF/YJUXZyzLaGk98BvB/25GhJf5Z1EKm0RpM/Yc5s9UawTiaNxq
dRAYkMLxzRvcSQfgqeurlA7/nIYSiZ7vhHVPLKoEGcwx1aoSQqOg6OWlJpC9yAJIfSJeby9TDDwK
F0pDbaOP8m4jbIjvkYUVvKKAKpaxX9TCw6yspcLu0NiC8Lko81fIvKU3PNpSC7rBPhFhB2Si5YTp
Q8uHcNpHsbXIX1mMTg1l7Z95m/dVGQb5cNhUwx6VmZhZp/2BnQLj3iU6FcwN/oi63f7rDH6sqq1O
m1tRUMsSkXXcWJquad1iEvarq+96Jq1UZFQPSv2BzGrxkzVFocNPdHnVizlZwygWXZBajo6GdqQy
caYkUPuphifGFxOni0PPLMeu6F/73o1ugGNssrhStuuQSKo9JvQ9y57lJOoxqdWf3mJ1WVaTJSFD
m0Bpu6m7NYxplcqcJDdsjby6fQmLHEDiOqv7mX6eoKCvXSdhcJqcQw+/sw6pQ7FOkWY7DGZ35yJ6
IoZ8StG7MXiVaZ1LDBxJCDct2Vy4UkGFZphTpeV/CmHSSZGV6JAYEtnCsfKi8LrHh8DU1Jck5RC7
KZ2dVA+f0t7qYpg+SL9PKWILRAzKb0KcECtb7fEURgjNXeRu6YxpeY0sqDzXfXGBzoUdk0ZMgEGF
WdtuJqqHqNKz/tOsWd4RMt8tG6M3LQxW7wJlweXzpV9rhfnboY4XnquLrTWgQnqiS8XfKgpk8wXh
ltx91Y7ow/kWP1ntXKZFkx1KQY90BCjST33TYB1oCVZaZKIce9XQEiLE0YggFoJuHigho5Cn8mw/
RlU3rAO6FnS7H4r46wZQOmaLOLd67X2P8Z31DkrNibDyO/MW6uZxVdLOks1/bGQaQsJlKqfEPpR4
Kp4jIAzUNAyopUH9R0XRruxy6Xb/4uGDXzPrhzGW5p7sEuMr6m0gHjtrLp3hbKakGpAmz4ssB04X
mt4e/ugcv/yLSxb1TuzeZPKZl7aQAwUZVyFUDAt0z+KVeZUs+f8dO4Z/aM7qefzsPmcmXIz68T46
skLLQZ/u/hxQc6/h/n0EQci/6vrTlM+ZQ+0LvieU0g8KNpvCWl9UnNdHLaGvcydIuyAfEmVTyqxc
jpRfaxZvtyCUPior/yZIVHDOtLOLBJjB3ZSXcFnrYR4yXMMVTnnZrc50+Ri+Z65PtCg0RGhbtld0
Ev6L9xj/Wmxi2iREOjzMtlvSb+iO+tXOPLwLfmjWJN3/k99iSZbd5Vr7IIe+JR1wiAUTgXcC9ZSK
r4P4x+cIvdtV0Er0uXkvHKmzFFHEgTduGn/XyfIn4KavRtwcP+tGatKW2xTN+uIs3IOyPdCTFTMd
slHllIP6u1a0IPhDPh4O3pD1zmc6aDmyPOk4crLLVFq/xddZDx5PnxBibGbzxA6nSCA9o4KS4nD4
Von75bCqTNzkBmPWFYhwNV1xqX6j7/ud9DIqlACf5vWxcwPqGiGajvJkJCZrtnlLwcbSiSj/CqM6
T1IvPsKkCYWTEa4Wgbfb/7moVmIGlLWkdk2c80jRZE4s/YuvXdwGeIWqTtMWB5TCF/2erBvbCEq0
0RZbG/dwwwksZ3BOKmROjyHwD7gY5ltahczznzuLiSQKfX5BsdwaejhMpsbxtfLrcT0YHlMsEXTd
UMUhXAffeyYSEOqRqAECxUfZjppODr0nObWJZ/TsZhIsBuBBo21eAD8jpQ/8T5M/hqdAdehkGpgs
7QLcmHoIXLRZeoNPKCONcQn7fnkQKbztn833XkxE0clai97PjJ1e5kncYQPzb1EDTB1DybkBzG1Q
2BPImakljoMz3PSsX1bxR33/IBSeJtOAWig7KPnDFGL7IylXlrhmgmOc3JvrmbGemLhUZZqM0Ey5
pFqQo/iC2HWjDYM9Orva3U25J7jVujLQoQUsLoWMChkEJWFeVLXsJpUWUEmVM0B65PYOTGMGITkO
8QxYxlfKVMajHavjpDELlY1xrpE4S2/dx5tu7hu0T6MbN+lzhTy0qOrpbIMe3dY4Va+oG+nUJSbb
qK48WImCNqlnUZw2sB4z+mSAghM2E1oBt5DUUJMmdPc41tIGDE6ztDuSf2imh9JDZOn1XN1IhTym
oQHQAF3NIR8fW2nJDU2mLIGvG+MGIlp7rB0HOjU0A/Is6B7yLuVVshxSADoDyIoFkYrv644oqynK
9RGLPjkQdMfXdeVciDXS4MgxCzHF4CLq1yZmI5I4G30ghWN+17+W8HvUZ/B5KP1PQTCqIY50v1FN
U7mx/a+Tc5NlOYPHX0WsoCYE/pbBD45KM4yVy67foS9bbO5mPzt8ZPYBmizRHwAje4WXkKEGtIUC
wfFdSp9y1dusGie03l6KcFWyCMtUFrdWnaIJMHxH4WyMLxIN6NOZStLNyGiZqdZeyU5tWsqAgpnO
Nm3jFBuTyo0JEbKdOGkZ5T1DpDwRH0TXwmtkkpN6quUhOagdSncv7lT2zky35xdbjF11X8o6bAHu
REtJ4R10SRgYb+0jweJRFgldYBpfqPvR26tlHOIWgfJs+43xU+T5U8iWja61vTNpeuuFD1dQio3l
a34nMNwJwvGH87+fpkahq55+n/nIo5MsO51oW1nJAjf07i6W7X8FOjtdOPWbXiGiHzsWk7MFAvGO
RoCWr9JpJ6UCk6Joekega5ykNnijbFfYjJh+iZ4DLEgwd/ayTTroC9Os05ONTkQurE9P41h7qpop
Etw2R/CNtAuKN9rf2/OEnf1pYdSLfQh2sNUyAILPiLCdHRtY+b6Y3Q/gBbcI+yEB+NfTEF7amK8X
dIiVgw7gDd528wqStPHNsNqF74wbomTHrm8xKEpl+RWO42Nb5xpvkRHOVK1wSUYayU+0ito+0Ps9
ETqh6bueBlGVNnhq/rLuiPU+n349IZdCDBubq9G/bUX0TDz3/qcNonUY0l/7vyjGQEc1M046Maej
P8mhscYjI04//Wvnh0dnsBtUzOKOwWzkSumlgC7YjXOuSGq68/Q0zmOccbnPK5+SN918fLyIb9jd
nSgogsiHeo8dkzx2RWvsl347yKoBMz4DYyK19tDqPMVvhSoGF1nvflHUaExWaytxkzwl1DuvBSDK
8E9UvBbA9V5Q61FCLlLLA5CcnwUu7eoRugiFe3fP+U9ZgUI2LrjO+bUGKc8KIWErCwjV1k/tZe8M
PABi/BroajbnmS3BQiMuF4QQ9rLpRmqhcPyJeGopLJsdbRjjeG+4v4WO38QqbG0ugIdcaV6NSJAO
0SqLn59w7sK5deTeAehAILdytWr8VaMKuR2AuWQIxKSJpTW+qvemID1wfHqqokRSAgUFXAh1Lyxp
VT1yPnRNUwyKLxmQA210zynNdYj9VJ5FEIHk7zWx4YLtNGv5/OjDj4PNyYLRrcDoPvA40KG+5q1x
b03kR2enKbHb2OMYEm6IlGpXQxgo5cDiirLwfkw1mb4P3RyHe1UQUhT8svRVjYqwStdvqwyL4QkY
snonAwUp83iobQehOj/MnL2K7MoKwQ93iv9qv4LjYUOAGMEcbMY3kY/GH+D03qc8rtrImLTk+2sU
FfDx99JZ25Toh+J5LnCqTHTe2kuYnqxJDHl9awWdIq6iBJEt28pmUrtaOy4qZHHeUuekXG5Q1UvJ
4kJ3go+01GuSImD3p0psre2x/6VBBDWHihJceqNgEN35YAOeJ+FbcjOPyMGcw9ZDk0774GlDYTbb
ILejDArZJlvvpy91zIz83X1/wFHPuW5R+82dZFk0aw+K5KXDc6CmT3jhAR63lbfjJP5AKQ9T/R8I
hRbeTkx7Y41JeNsmvoedd8zO0LBtkD3leLsbqNz9Jr+fhKTgtI10rcY+z6CV0sHTN9rZXMSMInca
0mXut2PZO4zlL5awfiU1PR6m+8rxqReM32ea1WXLelqvnSt9tnxd3YdA7LC8Kz3R2e1aOc07pBGk
9VcTr1cjdzEc0W1lDCVGxpMIUDsMwYbIbOn4otE57H8SmlM/chbWzmF8HSHBhEcnegTFhE1c638D
YA1K2YVbHbQQbRYazcDlp2MFmDhKD4XzZiHsT0E75foPfvOgvuJTYorzf3JmymR42LqWB2CVUvl7
DFs1N+Oc97WtMIXNtgkmmARdj6lpk6z0h+b7iC6cjCrmr73cPG9K2jtTqrJjbLEb3qoZspH5Nu1b
fcdKI8t4J6LV9XpJS2KBWb51dDUIE6eW4cxb1eEEXFOaGjAfGq3EoSHApUcEr206DLAdUMBDxt2j
FED/ah7P1RHNg6g/O1yq7n3Oa7MjnlL4CRUeULU4PtafCql6bG74qRqZp9Js7wirxr7+JZ9cZ5Gi
88BYs78I8vggS2kxiNigI7IEVl22XwY9bwvS+CcRNLk6AfNJmOCYnT4YOTDX7rP9RF7uD6v5EbQ7
ao2tZH9vUrhmsvwnb5p+gqEL/8gQ3Oh7qR0ozEccCpGkCOklcOwrGbxBpltl03L8V/5Lr7Jj1gN1
dvOd4FT5MV6pGKARrf4SaJ+SLO53dGgdF9yVcLljjUDSkdMOch+1CDqm9j8pFyjNkhvgd78j4nkk
KP9yICoutfeycUlzDdERmVW44MWPz9pqGrWeuGghOnxywi9vRDyiI0ZzPguOV2eyiMEcqdzmzrRt
0GL3zW0PbJrqD/Zj7fiefY1cZ2hxzB95xC37e0kd0sWrbc4U4nTITENWiiLUQ7SQRRcHm4kcdarn
kVf2GZ5oGFot0kAycses9HsbrAhr5eIVCrDICfrV4Kr33EXYbBMKkXFBpY76JiCadhiNMpTu0Tan
2utUKQAAeFqDmZcRD6mOqIrhjFh6s2CToKKL+M5qPbmTTFdYQHzCflcaKBpgODvQmaA4dd4j4f/0
+84aX5LW8pgJDE3UEdqWeK7m43KIeUbhUc1ItgPrxVO6A4au6AkBuAR3fG6pOCuOgeMNBLjRXAb1
slUpMha8ToxbG6t5eUD44yCsWy3qy5tRfGqutXYvX387KXYkzj88rQybMY3Xy5JGfAz25961+I1R
UFyRCGIGZtFDcCBw9fHxZ/uyFKP9gIai8oCSTi1NOUoCTX5EJPdtIJK1BwSK4UfhxhDqF8f2hszb
JK9NXYWVh7TM5VoJQHizNvpQ4eBSK9ZYERXVrr//obv8JYRPdTScQwHt2o0uxjRjbxuBuCMv1JHX
uLsSHWnHfLDe+agzlyQ29Hrz0EpotCpaZmvRE6sVPZJ8UOXrHQP8ZRKFvGRzpR0Y19BXZneYkVvw
BI1uo7PjiDZz+bET8ud7vQZY2PNVnsaQSlcbsB447a+loLLmsAVkIFNLUyLNKkdoureKZmDC1Q2O
3orkWKS0VjEZfKv9jzixbEAyoEXylp/TX+PcviysNfoZPgUCUWb+Vcf6sD0QPo+wkdlGDcCPBHlR
QHCZrQz7jRzWaRjF5x8zPMWOkUE8ctXrAGgWGC07ZeaXv71vNfR1bfNjoIVkqP5EdA6dyhscg9vd
V8g+RuBONsqOURTWRRzjWxGFCCLoDw15/Qtr1rEsgPFv5uQko89sY0Q/JOzx5a1gM86iR4YhmOb1
gj6Km1GAPFoZh4yIOcfOhhOvhjxwoUGljOslIk9fVmogzfCPwBTKqZoa8HbaNK3qIA436aqMGArh
b2Chjs4KB9tlFKUZGi0147KUILK5+gsktTLttC/8YQNszXLheQMjBflOUyGRjQ926pw1RUYkchOr
+2qAk9CPKfggv3kquykYW5fF+yMHKFLEkk2Q7JEB3DK2L36PXgMVg58jX5/zK6P4YXY9ytDtaGPt
38im6qyBuOMXKnXbXIDUQ5YiEyk95Luqxa1cvSgT53ZJUHmhE7NbeJYvuNUCmWM1Ca1NSEJ9qONQ
TUhyoCOO5gOJNtsDNd1mvxwcHxsVmJ85nQpmWNY8gn7ji3LJ3aPrijOSgZ0DtcsmfTJPj56HMtzX
c+Q+XsZqwIaqLO73fyCO27EYwpzxYBN7NqDO80OltzpHfLofD95k9IYVVuv7u3dVodgh7KdTEyhM
aKwiC8txAjj7QHa1Ckk4ut7a4YTSgtZGzaMNv5Kiat+LiGGnGn7IBhkd/YABHrFpSrXCKCLPPrlU
1rrcKzStgZSxEtOKLDecAo1U3g6mSrS2NYGytdUBFCICJ4H0OeBewYjYM33Rdv4imr+lDGPLDMXL
lLkpImqe33CJJfDgiUV6coVDxqUPzQrgd6L/NhaW7OUASHqXeAee7xLLY9h8tBL8a1CoVSEKeygA
uHpykRvZIjf1dpehy/NlxAVmIr9xJBsNuqglF24OpbUhBs7zTQ+OlIVHCQRoCCykO5HJ0Gmsk9ty
79tybbsb/+18o1vCTnodFIbFgr9KHn4Rq9B1D2XpXBW76rAXjo8YxH7aRH4/YcoMNV03GuEOaOrK
cRKg1hMG+MaDgRlzs2Dz1uWrhp8fedCY2EJ3RcTq9dPvGm/p35trQC4/Zb4YLIesarEman2UgF27
ZJ0+vyj8mrBpnLkBu6auwT4lShAIpZpLZdNkpg+B+bB8aigddQZY23CcFzRjwgmA82NGhhW2UAcC
u1LeR9346yoYpTR2irJrXhvNxdzbs64HVgf9/T2xljYWrQpviyLSItxReDj+Q0O8jlrHO2XQeqYI
a9m5pMAexinkcnzW7zJDvCaprg5c7uv38OqNq1J7afHXm5eecxmKh0zs5S6UAi4erAA577htF4Wj
zyn/rVc3GOwTK7RGoWGZWMy61lYawxoX9NSm0AcZ5lDm1wL/OGFK6tMLPqAJ2iTUQz7Qx9oLAftb
L2peGKJGpbW+jyjSyjXbBWegGMzJHy+Pqp1XLQpjHSdg2kTCFZn+RiB5NPlJIVKtr7imZlF/WmXQ
URvtpMQcG2dXxO/zhMK7MBjGbc/7LY/sxKqskMeZtFnfh7d1UvDv6RVbA+iVGzOvYoHCwH37zBLQ
MAke4ZF/htRYlYtgRTBc6tMr0WXyl/ko28gy+jsB7uxQVChd3Co0JZ1Q/LlpotfpSR/K1bklopAx
QBWOOMUzKAZGtIT4itv4RM+g+YZfjEm0k2rQ3NnK46QadyNb90fiKQVNS0HUKygHGtPdGU/7LXtG
3yah5zxBT4Ms0EXMJgLcfgsduylskoZdrwF/c16KBkLpF38yLpkjgVmRHYA1arP+1CRXKFKFOFye
8RcakPdey28aocfJYsxmuHs5m/2ZAB/Ftm9UPfIPnM2CT7qsFqGd5AWF2FT52boTDh1ydCX2mXNx
DT90TyOpkrotxFhJ33oSXcssqrzNYJtJPOxV183vjgbCVoSi7pSBwFfga03fqVuNFDMs2H+WT2EI
38v3/dDBh4R7NVTj4nSDT1A920UEewF6A0x+64wXpivxLE+QIdyOHBqVyhSX5aATtSoSQj3m7AnK
PbFgpRIpwolg4eqR5gcULBMftXt/oJF5l+oMqt0mwpnvYu2FVy/o7P8ksbll4s5S8GF5FG9RWnH8
aziclrfNI0P0I6mnA/b2SR1gZvQY1kgtsDp3gfEg1jhEQdeXfcWKRF1sgQLXR6Jy5KtXNDuMzQnp
rOMdQI3OspKzX4FlnmlZ9U235WYfbMF6n8Lo7iv/SonWrhx6ItbfoE/fJwUKDw/MtLvVDIIgDiEo
df/d7XDspjZsB9gjJKrLLyTgAxS9qRSmzbjZCNWPjPHOWTkH91P1dVYoAqPCUDcDedz/UMSodDZM
q/s3GJwPOadnBqtOUCx7n34G8FlHzNjPW3Ys1p0dFPkdsfa++LZ2DdLi15sVdIMBuwfHlZP2rmCR
VkofguAdImsagY82QaCiga3fobbRT8BunbZyVHlnesHoK7Wyzr7POUKCErrPQuqSwmuLhEdm9rIi
7RLK5iaSB4DWqgepFTkCxYg88Lelqdh1TEfEsU/R0pu2L1JObmVlyIp88HBFbGjWPEvO9kjMAZct
K5ZD19XuHx7o3DnGX9ayYU6g01aCWiRYqC31P8UREKWkqTbwD5TV3YkVfvfgia8n2aOLE5pX1mfH
h7erWUcf+UUgh/I3HFkawiMx8DzmzJI9HjfSDUi9bs4bItURj+nEEqEw3pgMgxg5aznXYEHjDJN8
7jRpKXxsjB6y5fyWjjRuHaiMNi+DZt2wEXJ4ZoeYhS0kjfpZ2jRwi14hR18U5ANs1gihECmCD5u+
z+3VDG72vhFzmlkmCeUQtMCACfkM/lDEJsjnX+n/41+lhOuwvwG1eJyg1LWrp/jSroOskNQDZb4U
EYZmK3lblk98CdnL/jMKX2dAeLA00T7eJVfHbhLlklaadZcRGNzAgIAjXbrzHhXuBi0EDDc5RXE9
eY1DuTxSbjzQ0dH0d2oJfXf4mKnvYnf4xNbKPZrlsanuesfrUItkGTRXFotJpZkoTbaoytFjQSX5
EJ5Agbgl+ZkhvCSibL2DFyIto2958e4iq1srJIfxhwE33qkhK8RjOBv5pVoVrOXZGYFWHqlB8aol
1j/nrtI2w2vVhQmH+w2/iMJ+OB/JfVwhTKXUEFbTZ4xWG9853EVrkTH1+EHit0Brr7jQc0qAAzE9
wS+gq/IDEGGqOR3IqJbMEGz2PIkp0t0o0EGTh3uBxR4csTwGkV2K4GA0IEHunuWCUw2FaSY/iKHd
9oMyaNRVdO8Xq1v/IDUsgxktHvwShi9r4QWaerjrGYT2F0vPDoG+1jTvMEzrj3r5JCKSqefgHmqO
mIHTLtF+G7ha7GqCNXtwX6cTCjr8u35jrZv9bnmxfmpyg8npBPMEu2fnPRz29PVsJ12WYR92n53i
uZW7Zup5bjv2FE0WSpHNYc3cajQGQ9cb3t3NYiWep0Xl8V4igAbTYvE+KZBzZLs4DJkCVBn/8EiI
FWa5em1TUZQ43msoBKP+JpPxE7DoNQPhfESwX09bHimqHkuCKOxv6UGm0T+PRko2dvPqbbt5rRx3
kaL52SnJUmxFmmsgX/ZfQcuTPvx2mVqq8Zr34jmPxck1BTSX4n5Gb6TC6uGJJMX32K5eFA5HYpXX
E1eSHr40YND2/w4eFPuIVDjDsanUVPPWbfXvT3cplyqs/92dru81sFe4cpFeFmy8TF4PX/D4rvLL
Uf1KJ5S6b0amsEPGh/gYEdahNURDIjNaBlWTGm1hgkKTY5ir9azU1XzTwwJ1snbVgDhIQUV34IEp
MTrELEe3Hf9UqiNiXGVQFwci9zW9LyJiEP3r9Jx9WHXbO1Kq6Q5DatTeP8podxNDidMYSbhmEw/2
u6Edcx5FkEBtWqVd6DyzVnlFYj2JA2HigFUiWfKn7d85WYUik96I8PNuKEL4pqOiQpxlD9oIeV9x
28YhH74W2TQ4i5Eku5JQRE8ZonYQVH4woaXJK4CE0YprTZEa+T2qi0UQ8PaoJATTqD18n3k8MUpT
ioDmPe9aLdHO6Cfah2x1PUXFMni+AYk9iPDNgAtbQf63RUVD8KWPYSJ3baGI4RqM7bG3sfInhZu0
vJRBBHAY2UsaUW7zl6u0KZNt1sWNS9NZ/1IuTt/jaA949x76PIC+M2tT0GZpcvdXWQw5S/FnB/uL
C6U1GJRBc6NYWAB2oGXz1hYWzZ9rDTu+46M6GMDfI8XfCVP0ozwJqjz1t1P7inSceCFN3pPUEWTr
byAqayNLOFZiRAfusBH19pe4j0X/yJ7/MeQtOulw5uWK8DLWsE4AsicMHgF6DGOs83iRb7TWRn9m
Oo0XOgJ94eQ/RBaCSwtokT0NaywdGMLGU97S6e42Y4Yb3+85PvM4TmfKfvcNlgnnUtZeT4+ecfja
DjkXU8u9xJ9A7zUO14W4hXSj4UOvXMwzhc4YSOrt7Mh4+vvDGvz9wdwbCaF1yN9odBvJjM51ajPO
mavPnpNsljQdMJ9VdJxgvRwbarkIt8xxgIfW37jyQWLRhZ3HYsprJi8EWS9FUZvxaT63JSF6xEz6
8xwG6mKxgETAmo0aiUceQZh66IT2X6seQBUQfRib7flQmGpAy7WppPEFjl+6ZmqMFTJ6NrejtnHk
A8b4Rlvue6jXrnMqT2ErwxV5jDlC71YJyPPrr0UI6sB6wmmPZfL7T9OkAn/fX5omYHDoOFKV5idQ
plwkHHqE4q3P3+Gi7upGyJmjOGSMyDK6Lqzgl4bXFx3oQ3Xbpi8ZivbSurrcAUSmHOzZ3mR3YLda
cxfFLDyp+kEEHLOCHYINzLQpsNmvAKBB3NB+pGcAfZ5PGjJDQa6oBMtfTBviAmntnpxTCwRbc+B/
ECUjHqTrMnoz5Lx6Cz8T+/sLK8MH7WTu4NrjH3qQSUxUlghShH4ygCQM3HYUAmq/qgs6KhOJ6Lt/
M0Ckf8lbQqJuPVYZL6A8iW+M6nJSAmpITo/kwS9ir30G1bV0i8mMlJ3nBgwXaqgx1aM6fSzy65jZ
nJLvcZuj+5vcmuyoHd5Jxpu0w2rEa2pmFFWI6a/rRMGtTNggQJt8xUhP4hI00IoLdEhtIYvYw0N9
hTS95iwrseH9ohpJEtLYaC8JZ0MrRMUlavEH4wP0AJbO5+n6ZzoETCZ4aol7E4sTH/Lu1nxrknbY
WH0JukX30R7hB7YIePeXIGDWuPckYV0bjbvXDV0IM7GY0diAH8cr7A8sij88RCTCoC5orrVc7JK7
tbaSf6OsqQK7XEr3O3s4zzvYFP2YY7LNmZeK3bBop46N8bgESfxKPlxupTmlvE8394Ao8ouUkS5o
a7TcXoqklAQUdY2xDD5I8195hZswVAa9h6HyOBKPtj7RN4AIBshPYWjLh3RR+VB0SKk30tiYl5gf
ZZUod3QfaE5hTLPIMasSH+7IP/eizHz4cpXS2AXXNjGtdzW1ZrmjhBCTwjeNjSWUTbNHPMQ5Jrw2
FaEe+FBlNCxZx7JFd4SSbssEifdjtaMI+E5SpOIlshM6jfpUPNRok13tDQ5wMU3v0akpeJfXZEXY
AWSUEdFzGMp1cAfE1uOYjDk0ONiz/8KYV312wbDBjRrqSySxnYTmMRwUD3y9FGL7rzqR3vGCcCPy
/V9HA8ECaz+dSodadD0vXx/zvfZUUPqs0TcAufcdOphH/esxcs4aHMGPTNKHueSoRny/0jN/2htx
phDWfsdD7pIOfka/cUGixsPMl5LJTlLhEu8SVTn0cn37apqIPUefKuiaqZdlEoiOBmAjChk3pAFz
MVdnbGkUqTV6rXyWt/FPWFTaUdxD3SePc1PbSiGS124ZWMGHlALuyvligiNQ8EYuODyNYOef8Yup
z+HoV2apzOCMU2F+OyCD8JiyyMEhhakxAW3lC5QmSFIX4315Y/zUmKWopXfQl/G5X2bNp1aeWBXG
tjf/xXGFtAb4b6gJwFHUy7X5vR5cXOXgbaN/vl5PzgDJMO087BqNVT/64DsNgU+13j+A3Cj6Bsma
/i4QjmNdpBd9Ij5IYnSimBATY16mGzbiYHT/tezQOF9QR54///DInmUlCesZJ+vh+pg11AnMKmRs
2YagtPJaeXcBpFS0J+UAxY5BJ/vkV8B/Ys7ng8VMWQOWLCYPupFj5FUZMSWEny7xQHKYn1iqDHzR
WQfB5hE14LOIjewXnJBPCK8YZRtOY0sPjclcAiegv0/5OV0N5VN/V85K9Op5VKr2LSDuW0tDxGl7
xBU/bnrz9eW6Jx6U6swm0E2f3yz8Kc4dSr1+qS+hNrFvitMv/riTetPewVU6MsMaEi7ub50u8KqQ
x+3u1RcpYTKUaOOjgMCkQbj7nh5nTn10eQqBZN52WqFyeFzn0/qU2PS9jcpJ05RJSm2gagR8MQB5
Hvdv4hwO27Ub985ffEic6/g3VdaScenYaEQ7K+Y2c1Y8j5CX392xK8BaIjnDFiQpEtDoqY80Rg0U
BMnPT0kQDawCCm/+89CmGngHYcpgW9OPB6qOwNDyquQttt124u4wYK9A5906Qp0QXk07duf9axsy
JXfzxcClmRvbaIDxInZjnwbeBKzeVhztlnT3OaxeIN5m0I8wytQFlNoCVhIjDpVMMGLuSLXiv9rI
XJU4GCtHs02dAwKw7dLRCrjgUYq9Gmd2m+WhOzcNl5mHGDAzodS/7Cz3s22vkw458KIfsxbGLhu1
001gmJMTpD5eIJYuyuscGQbLlrIIZE+YIhXNh271DnswY307DTzg8OqT+o4dxaEcRuEfsJKwKmr2
0p+Yehtq0rid42DqynVCWR+GfhtrCm0/NmpmskMWxid3O77XkSojBYiBFCkZZIVx3tzg/XgnpnZw
+ooNVAN+awOWefEGTWNcXD3RVeExeQShm4SseUEyJn4aVqovNwuHF1/++6t8x/uDBQpeHZnFYzR+
/bB4oYU9Db79TgKvVFkF2zk9ld2XXYtw59cNnGqbVqdUGD0+j9XF1xXolMsfZg9H31Ld2YTpCX6t
eZsUmEdzAc7aVV75O/ZAYN3+2jNRPW+4yHEX7TjinwCzg36JT58K8aSAARSR1OljETeM1LLhM1a3
ZRcihJ+wVfHs/Gqhi1g0Lkuys+weUzT0LubQ4PRdxjwc3lA//xbtSvwkIBHLGrQ4zmktihg6RCgH
uSTZUPisJ70LluDjzYvHSirEA9qrwhGVLkUUr4AsHTxycYCtYDbkhdecIE3sD8kYo1Mahs0yHcrK
x2pZBjMTareCzzqVrvKzYLzMUUMyNjTLEQ7Kh6n8FCmdHOOtyi3zCO0o2n0Mym/QZCcKzGclvzY6
9rVJNn4m4Vqa9izVB5I9X6Bw+7tmTLLvtZQnBa4MV7FQsauqzhuICw1ZssBrBqwrYuSrsTO96zYB
+zd8BQSPFJFuwWtoJI8i+teX516HRxoPqgezK3r/uiFyut25FOqg9+TcJ4aV7FjHsmplbo+zKmh7
KvrMNXKGFsN+61/11RdOT+EnwOGpjboTZSSQV9HJEg2mDjTLZuOWpJb2EFXf70LFtWytpbq7HR1j
OvbIOIrCdS9lRRHvsPh1A6iBisamwzNaU6s6Gibxb6G3LoOLvSfOIepv1O+IIHH9AG4UJls4ZkZ+
q10JcHL7byFxdW850/xWhLRUagg6I0Spq1iwmgFD0pbEWU9LbIpuhdE9pMDexXoWgdqJcNNd8JFB
jvcYc5Kv69VXnQUFj1wUo2qNfCLRkqNW6uV0rRd0s0eTKbbOMdToffFkcDpSGe4yw7hDGIfKuM8C
rSRcWisRIyDa0VrJpZU8sxl77J1mLSBsTaaYerEZvUk30UGHxHX7x5LmHVhEbd/jOQc4YREnx0CS
l+u7pMvyJMEcwV6goWlxtmTTlw7c34g9qD5vSjiEsSkrc9gOdpvXCW/6H1ajWxoGMgbEJY+1deRQ
zpUaxbXsYVNvwJjVPo5+I7Ya85a/6xR+ulYBWTEqbgHGyxZSaLKlGozIo9gddXvUiSD4vVbwm2HA
xJryYRt+lNW1SCiB7ghaHujorSxnZoq4isjwpRly7498jPy3KSNlRgEJrbz3ZwKKcHSv7oj6ApNx
VxQvRnIc5yB9pweVZA0kYS3/K0us6kjkTs/jAE58fZcVbQg3tvZcBbtHKeJOXGdl66IUXenwGMQ4
lufENo56GgEg3bW244I/YkwX4c+r6PReay15c5Y5IlvfNLPhlCnezB6qZRz3NUFKwYNlMwYayLG4
YmtEHu37mNGtIpm44Dpcldkj/naPNDpQLJOtQHwmB+k2VYdEmcDNe1kQY25LEQi8CIzYGYb5+xJJ
BIRPw3pn0EapzeawpMhZTVRDw8E4EfwncZSGlF4JZZYanaJW6PKqj9FIRwvzqJFMwGOaoEqIPUat
k0DlXHNQPlP1bdb50Lt+6Gl+9ZwjZj0swJ38BofxxPiMV3FiPHVnkCYXp2NLsRYEANak5jGXVBc9
D62Or+cefeZScV2uKQfGxSnakc8T72JYQqNjW0dbuM8fhjJiTMa0/HDCxbybjeXX4SEJSECpqQ6T
xJMTSkZ62sX26jsT9gTxftSs46/LtydABnFxkmbaqg8vgtdhaMA3H4zSPdGv240suq8i8TAzIjFp
mjHLNc6NtiAQzOABT/ot7ct2g2mJcV79uCPhXjYRxXS55PWYTfJhIOhmkKtp/gR4mzvwswCQZZDk
37MtPGYSHifqEALXm3dpqmcd/n7jeO+Zrhf9TL61xJBlsRnVUf2uMBLT40QJmDahs6QMqKOvWshY
8CWnEJv3Ca5IgB2JmqndsdzLl66JGpepn7Gucw7ljbborrvGjk6N0GAthYcVlkZF9ZBD+8NHdic8
c0yrGp5NqAf7eZWVf8LEfg8mEbkkmiq3bR1Cg3KpNwheY7ydLo5jNN9use2tmFh1/++D9AWlwtTf
PRekKT5N/d46OEVehHEb+JxNQ5Anzf/CaTnWFCIaOuytOmW1hPI/hMx1GlAC1zIFmgHnxugIJxUk
J18s6ilEQFdyqjuXCyCumy3BJ8Npvm3ewfgbMN313RtOUIaL+UpmoOIFXw77whBSMpUVRpVB4FNQ
uVnV2y5lVDMapfdv6/bpobvNawtoPu1bDayUI/tWSpZtRYO4foeo0pf00zUlC5tf0wQoItAm6TLz
EZ1Mja9LGQwvE3RsXW03wqaTxfpXgIbXC96w/T6c/ZdyuK/gVjot7uWp1rOQSnWFjLzdx5NLwCgG
Uiy3OpM1OsGXCgD7Ctf0MAbqQZ9A22YfkGlEd3f/VGsvZa8TZ+gb3ZBUMEnW+ZhMMWIQX/Pl+osh
2R4VlRcwQtSTT8fFBldp6a9ek+L1iayqoHv7X2pQLsM8gkl8mEQFT5yTGCyTT4I+AC9Qbwd7mMxU
0KV3YkirmHLPiTAhCrHNuxG1vWZq9yBwMBDvvhW2fYGAJ0UWRCpWjvbjn6z8tFVrCTFuFQ3SZYrF
3NlBM4rYQHoGXYLj0kJCSNmYcMvKHGSAtxYkYys007FAXwlMscJYpMu9Qlx2pySR0iiAVvK5r/o2
Pq2OB9ZRLthm2jBOHDfFXgj9SfGw3J/OfWK0nswp41uSv4cHeDyDcAZNGYjoBBxndhvmqcikjFdw
4wc3AL7at3WeyjTBX0YKjgqL89Bo0xBYT6ssaXikGC5nYK7ekUZ1p7k47gEQnmspyjy4KNEGKG0m
epx7PEFHSdR/aIuIE0Lbtg11buNNugKUmKaw/nzGbNv4ombi1K5klBoDqBwSZoKrMHmWdPUy+TQO
KLZ2N5bZXo1dukWuq7ECeJNeqtUh5lGCvIxg7A0GPHA5lcMfamRQmlYBAk7/cPBOL3k1qVrXrz1t
165t1wa6zXl/N8j+GgL7VfIQk5s4K6TH7bhPAv4KrVQ1QTbdGCo87xTKLRAT1rJedFny/hq5nDWm
lUd5Qje51xZ+BNM7tI63u2HDWDKLb+piRVgPhcfj0cdOjXkmcs4pFBquzTpDN2m6+qGXji4T7b+R
qGOgbSOC8EGxs77ZSTSz7Ba+FXJp1bCru5xlxRHDvSaVzDp/6M3PrUzf/RG+rU8AA/KjgqStQRwa
jnawftYYxQAvtrOc56QEcyf6NABmvTgH48RdgahuzkehBs1WZQw/UKn8QSE/DvQBZOhN1MkgfJUg
kLaUXykTyKtaECnV17TvoNZLR+9iTYEulJJdRosZtVhilf8RT6+O4BingGn4zqWYxSVQiDp9jufT
eG9KiAogYehEjRHM/p7U3gwVKegWdYdIgKzGKsEJgE1NbU6yAWCf8fFGdfsVvnQL4Oo2JCjl/Ezb
il5DfAkenc0mhI3XvC1howgZDAzU43eT94kl8bg/lygmyTVZPEoJORmVm0uemURGkZMXRXpQGdZN
n0gstlXlt9k29boordoKPX7xSPJy3swp1i72MwQGK0zUea+Evp8vdH7b1VlU1OaN0gYErMbLMfMF
TOb6r1BHY7WeMIRYkixUP0O3yRcNBGjEQ6UewMimjzU/tUNzyToJ+csbLgdVBYbcNNtpyR4++2N/
eoA3O3Mcx29YL+P2K0O3oPwK2af01vc7zbMpfhxJGH/dgpDfd4kdCEA+btTjYEo7DL9UEpj4mpVA
/tRxRwq78Okh9EK8cS46XrycSccyLb6a+3SrOXbAouGjHncEKSXcIgl8frAoogDaueJBy1KeONvK
h9js4B+qsptVsAh42r7pCFOn0lIIBZDW84/K09NJvkClF9F0XQyvfMzL6CU8ECfFD1NjguFc1+I+
mPjqgbPlxg9DgQUR9d+LgTaNLoWKmQLglZU/gwvEBEL7D0L2QksWORIdKlLR9VyA0YkVzRwDMWVb
hn23ZQu8nVvkMqWMqmVANuYVVn74BRFq4pJzKK9zK9Vc/oHXLXVYu75a3R6MSgUs1bCZ7J/+HZBf
NcSd7AXPB/95VmnQI/aFhdhg0fc8fEfoTq5EcpKtseeI9nrcyd/4C6SnzfgbLklAXEVS3CCHzybW
0dSrS+NTi8rH3Qz3J+P6pkVPyDWb+5kO75BU6JIeijNuQwsOi/5IrFMBjRuX8kqyMVVknYIsWM2N
CU6OG335MWNykTsDHualeGFMaM+xgBLKdv3QgUHhzRciZcIUBvFmHcCOEDFAQO4FuRVQ9dCz/55n
N1lFodOQTewTqLJQnfG3xKJITGIaHSHxi40cWIoiuXyHdXcaKv9D/cU01nSCzuIpXhmxuLCUqP5j
zUMSLXobupt2Mw3qibHuwRa7Ew6380cC7KpirOVry75cqsQL0K2BKOCZp4JvzJkTmTZkaiUQHo1L
3NO2J+/+GHBkThEKKpUn7+JW6XKxnMJALFV3WUqzT/h+cAkYeZ9c+F6nXPUoQGy+A3fi1U4rhrQM
KPT1xcuY4XUVQ/5vj0lrXvLs+u1ZtQWD/R1GQ1t0FwnrXPeh6KP8Ck28AGtVHyx3nRv2D3cuyv7O
NXbuu5J2nDRWU2LIucvLJJqnqRX2iv8lTXKZ8Jxch3gsEDerf9cJ6nhZHzQ8GANYXPiOk0B+YhJm
9eecHIc4OO44KYJAY1jWsEAj4UbOyNXYYXU3qmQDkr8IoNODRhw7I6x3Sh/NZS+8AjcHUMjtehWm
AHau51rIlAAFax2hq5f/1oZ+aqd4mtiw+/oMfuRmeSQSltRLeeyZvfIgk20j8W2Ups6d7WOMFZGi
c5mY2wxRFYBwB0UGTvWqOvRi0VYxlr7NSLH0K2xHfeU2D0QgPRIjDjsLlH0rrN0lw+JeFSfpKYr+
k4kvJcDIbqunHTlrQnDBkYv33kW/s0TU/chi8Dte9YSqOPOhL4BwHEc+8eNiGsET0wOM9k6tRKYA
JdZ5geOb2ppu4S6xqu02gpPIwu4Cj/eebytUbTk8C/dRjwyPVa18Hq461Ye/ZJGmI9sMPJSw5Itt
+UO+qieOyvlxpwe+TWo5Maa1NzvTF4ZqzXW1RV/4VY4QQkF2136A80CFWOvJpE/Mr8yHadMPigDP
2D+dID9CBcjE4wLQyJrQDKNOTfDdme6zcJEk8QuX3WgVB478Uep2rYa/fhTTZU4/FVsO+Glsv/XR
9spkaZ+Y/2pCGokL+6/lHh3U+0gdkFky3XTd4Ss+huaHpsX88GliQe6u7KpVuHKvCiuGxFKyC5Un
ya+JKuv0qjnZb82UVkZp1VJBPgMmIFDAzio9nFu0Fx5TMduBmZgjVsPAt0pIkXTS0syhchB9LkcI
I7pCLNP5xV9lWeBsY++Uv9IO6KOU9gs2yUfSQtMfnLKn3eAzUf4zu6+YF1epU0dl/TIDyuF2a5Xo
XtTvKs92UGYxOjlu6VwoAyrTydUxg6udW1gV3G4989hUYEJgeURYQwMJht4xmdxYWtSbKt8f2KkC
13+5K7EVrGJK2leVrJLuSwcdsLseKyoCOYWrFE7bC3UhZea5XPndCcS5xmL3NUbiFwddAiiz5Xho
sCe7TFlq5SS4b2NzLoMTNXBB97EAun1ZGUWxf7L0RVrKHPyKJtEkwaVeNLaHl306DymGw2zsvf8J
onPUGqKREwuY/4ApzrHpCI0wskxRFYU+vLBEQbPjxE1rjrV1zwXRj7HIHcsSrHK5lFjhUlzqyNY4
DUqr8rrKdMUjmRfckGFX25FweJTJ3sabAe129G4ZWEIqLCl+xIN9PLngrIz1Eq5bQqFrlvjmLv5e
rL+7SP7qWBsZOoCs+dv2z4B+jT1WNjF/wsYi9UcBP37z+ZAkVklC8lIe8iMpzP4sLQBTy1psj+aZ
grsnNvD7VQRkkE1mLOSg0vI2B32NbluJH5PDJfzoYtBBlxifj6Yr3kSYbVealMTr6y+MayC/0dH9
6g4Jw2ovvoVzysYRbEQ46NSXRXuVup25Z7IV+SL8huNBZ0oG5PkIWbq+iQd7Jwy9Tu7E8rCUnQiI
rmgprwAkfrls//OmXUGW7zT6LVRWxYwAegTrhIHHzc2qxdMQ2rp5hHODrbkAtSQLZmUQ4tcZRf5t
qj0BtqoTPyINTiKmLgadGvOF6BmQoc4am4HmGlGffNnzdHdX7WZgW4Ds9AE5vB4ytknbPlP8G2GV
VKXsfR9n2FrooCqQ97AFwOw7A9nyb1wLq+k2ce1tokrqcDm9HG78KL6OCzIjELNXLb0NSD7o76SS
gb5F8eG2kc5KzxCBZsI/Ri+kNvCGjBB+84CwEYK+7YJg9bEr1pfmDj2oXFO58nOKwLY0ARJUA0Zr
F4p2xZlmYHQTFM2vNIZTaVmie6YW0ZotJYdC7xytEL60XZLZ7R2qeOxF0DwCnXhjN0uKvxd/qKdG
JgUBknqUtBiGtAAxWMYzOxEQM/k5fz/2Su5ojrsnEttt/gl11AHnvhgasHabzp1FnZl4uemwcE8G
4uv4SzE+LPVOXn+WdbdarGOLx1j/r9Wxdclk1SCrLmW/i32eutRCEy1VXGdpqbEIF77FZ21Gq2TH
UqxmaJIoI1e9d2803wWQttL2K9ceuZ3zfoIpH/aH91/K2/AguOVJ7anXqznMkFhEn1THkg6aY9Pw
Y+yRb8nvaZjRaYfTqsgtg1gVX55td3opYa3BGcSf6+JGdiqJ335F7MdcatO4AXiSTL38IQloEqwc
MXGrqEtpTgk4YmzLNCxD8DN6rPvvtiI3FWsnEJlNdlIsEENsr3hZWAb9YsrIGk6oXYzaCkDYUVrb
QRBKvRMadUwlLAFC6+3ovPPbsOO95hd6KLIG7iq36vy1yDZcVoyhHpXNzTJWO11cAmLBhthiJi5j
gst3eBGHUMRx7atjPJbBkGcFDosSSmFTQN0ZN1yufiI7fJRpitpy7JBMWcgKOIYhN8asKiXwdSLu
tNoJtZyH3J13+90kgbogeUrnSwhMn7GFvlCvKEKFtihXdMuyTerSSRM5qaeC1P7U2EZVwjOfjAVD
e4uxDUQEeF3o592sErwXVgzCueL8Ci67TVXEgUNx+3zwjbrhYcTdLfI7z1e6NLKdFvs0PY5nGVJ6
lpxCsR+fXqnlVyYlTv4PRo7NEA4E4gRbtd4vlonxz3DIsFrxm8SZ2d1z+6zLmeOopggzZ3qJ9LfU
q/zekGYPf7x7iTmEjFgd9IAyMSmFMTLv7B4xxWVDGjjAZbrbAz603sLRMXs3ePp8BkBscldOux1S
Hqz9KutqFa+X04wL8gAg7ud8WIYV1EJgFOZXflNEINKCYcJO2yHQbYySdVVICAzrcHdjQ4yjtFNR
K3oiNAat+6q3eyOZ04u4GV8QgDCax4X2JJIDcJRDwllOmaW/mAMKtut/wsUe5jBiT7g38LGCKoXD
GXBJvEVxNiTHF/hVZhhpakEWZH45tVQsSKFMdZ98ZUzpOUGH66mYMAh95afWkaP7sBve+t6Wr29B
TFEHJ/mJmWh+eYdUnxziwuByKRHUxNfVYn7164q8H7HP+cGS8TQE1l0qByycNi7q/9MRAWMRel6q
K4ugSqDJCfSz8OuyaiUDcomB7VMZl3OifG+0W9Joj5nOqU09KJPGxZxFHwex+fHOwZYIjZqIOPkK
4j0Ec2UQATkjtr7WvUvsQEZ7I5qjJUErg3eE3ceOJ0ErvD/0/fadFZ05EpuvbDfhCZzGOm6hPZ15
PI0gJjxz7y4GbVS91nwqBAKU1uXmQgQC25q48WdcV/uJdfGCSrUb4TYQ5UuPPRpB64g//9LdNYMZ
h2zzq5+Hqq+D6bI+GzArHPmdTSBgGqOe8Qq1w7PmU2CTkWFbqQ/BN73UA9gcOrAAMNXPtPggla0+
gAz45gO7jP81RqQF0weqhLMZAmqKQQrLv9vPN7oraB8/J9B49k6Z9/QqjqyyKFJauGSETkDMbTtT
aDrPNnMD29xXu1oWG0zGV8JjbpUmcjCgTVhtvOrrPj4fOS35Efpa/WVY3pfOvvU25HCVeuOclDl5
PSU2dTrdjK50VAhzmwbLDGEBbQIWlyKl+/0/yVox/dom5lGsfzztBcIJuKf2xjY9LGjSafPjnUpE
fE6zzMbvycTbDMZ0v+hoHLFTJ989H3GAwHt2rWkC6mf5ZlNKRlnMucdZYgTHMxM+BdQsZ96RRNLF
Utdgx2egUPjVGlUbJFsIohw2DEDjnKdWDtIBBA13JZJpvwWucdBpuWPnTKtfqXmxz70xs6wxAsYg
yb8H5AZq/uhohqKBUCNHiabaF+6ND297vyXPRh2dP79het5FST5CVlwEAZ5ORZ7IYD/6+CfNj45T
AkSqbXSRqT4XuQtageAeUA4YM/vEBnrP32ZmlIyN1+G4uWIPM+zhQ/NsLxejNkT9BQvv8AIMM0u/
JXGVVbJ+9zavEnccYvK9heIrew2GviS15ZAWSBGO3OIjIFCLaCKftZGvFSKLiTJKEyEXLUfhHI6v
Dur7IpgdpyniKV1eO7zBXJBQbqVRC++pm+pgRmIzeke7QTtv2Du/txM9CRGTXRxM/T47Ld5g3oBW
X2GHa+oqZMEAZ8FrpJoloPdA8hE5AvrLwBfyf/Ys82/8KcmHCARkuBsB1pknbvNxf2AfyRXpjzvD
ZqRaDH4afTngdRYvDYhhuCHJGI6xGsq4sOOAd3rGyjDu1s7QWpS1ZglxV1SurIkPT9tkzBXhaqiD
+XcLcB1xih+z1fj1+k82GHXm3ECORH1PNWLNQz2KeQjM1Rr6Oxmx8mpncyvrHdUWQXzPYXt0qVB9
DV3DuE5duyL8q7+Ch4tpB+YghMVbt7pHgJdTWQnCu+Snc1hR7KXEmpV/giADQidAY+7CRcymJJyf
qyY9t4YzkT79ISRfuubYcd6w/xm29K987hVV4IZO50r9ahmiZdBnoA7R0dhzvL/pCYFpPPaB6huZ
+Phl9gIDQ7t9iedHCem5PJhpk7n858/1iF9c9KR9WFUwkZnaL/EJPja4vRM1cfksmQhYxGkmGzv2
PLsjvmtxmEFB2DzoyRtiHRwkJ767m1ZxLqaG2PvwslcHV9ev2uCteng96xYZLdW+QNge4eLWA8s5
OS3w395mKit5gBr/3L8KchZwsQPV20S93PB0icMM0ZB3/QmkQ4naFikTVi9LtYKOyrp2mGF7LMj+
Oe4LRIAVZ2QcwwsJC50F4cWoxgz8HNIe5uAOat7W1pKpX7Ykl3aWqTfo4rrbqfQh2tVV5lWSNUVq
WR+DvJunmU51FcO55EVU2Q/RQekiQglTli49z7lDT8eq2+u8CX60ql2gBsjUxP4toGx75dHhX44R
uDqPmgPUWbFtTp/WhcvbTTazHWWCwS9f87yxfygCj4cdjfMOiVx0gCoLny5f05TglhlU6Qr7gLO5
nRgO6RmQx6XaUnjO8UBN+KeuxJ193/Wc+rMmLS0Pa4YRqSjHuzHKmho2bDFIumEv2WY1Ug+ci8MZ
45ktAy7dL1P14x4fsdhcln81bXaZA+yWoQ4UR4/mMCMCHrh66zsbh9lCpFrQF+w/u44/KWHVDxZ0
KsFwdpN1ePwzk1Ul6ZsumOV9ZD5Vc2yN61X49m7vQ3YVftAxq5l0hd5IA5RbGEjgUXxOXADhnU6e
WqxyzGN2pkrxamnG0MQlp5Z8mqV04jnzZ+/7wslzDC99xw+Ks+fu4e7RczjxbWP1vTxkx3lCPWWu
yCdUlIY1lrTqESWyipxSro4tbDuYo17oCcMFATy4OIYfGxqTze0cJxR2tY8Rz8o3CXynX2YxYoBx
wPLq+dMxP1yv/kU6YyPdmgz2faUXZLEEGxsib8XM6Ieh+6tUl0oiq1HXgQNM8Flw2MiqZ7vxHGlt
4HvnTm2PHCX+7jAnJpf9IpiwVtIWluLl/NsEXPNXbE/AdRDBRZDF9MWVKSb6TAWWH5ZvsvNU0n33
dLKVtZOaW73zhPuCJCw4TQd/rDHQ097hcMY83RGhO2Scs9uZ7vq7MhGmmFZn9QSIDsppoD8eCbW+
1UsescjzvmXRSp0rTGIbBpyRLlQm9I6SDNhLMtmVqbKpy5CP0PWpg8rUYUHulVsuu+7VOM0pcCtZ
I9Sv368ibJdAc9NYwpzAIvhlYdu2tqeuBZSyf0FEBh3m7G8bOgXUil1IgaGHDWJ87KU4qBFUueT/
QejIgH9AXitIlWj8bfEDkkDMOF9jweAW7hnj7wBYfug8LEUsT9AABjtVXhxlHIF3CLSfde5DIYPH
7qwwFZ3/q7W09uzwdOUimMOXVCe+HlyEAUi1vjbRd1w7OTuipWWYVnxMlqeruOoBO2OrWWVluit4
47dstd3sVYa/2d6jp92ysuxl5L/fg0gwAzMrhwsalLQrJsJODgMuawQ/D62sqBKc7IR8FI2wG0iV
uvMCaTfBLVdcFCagiMRPxWN3u4pM+zM+xKqq8TfVhPCt6KccGYipcdF29Of17FZaCXoYrz5YuURy
pTUP7fGWBv5hVZGE/ICo/TP9FaEmTXHQEEP6oNlx/ZhltKJk7Rp6wYBdO8Vg/gWelt9NBGPtN5Iy
P4heCTC9fcR90P12Rx6T8R5i1DwijX6i6WeUOV7TmpWwozPVJhfINLJDEliH5W6WWY4XpCTanpMR
BpT5Y4pTSlPmbKH5gIUuAuEpwrm1Bbv+h57vxbMKEHWBaYBUTQW2WG+L70kfFRjh3p9sPavVyAsT
1f2t4eLTj6QlnhSlVWcrHfhOU0V9Yw9lm6qq15sz1WMKXUvq0AxOUmk/+QzTUSHYbtZfUX4UY35m
faGkJTW/bt98RThdNh7VaBxDZlYzGmHDnMPd4nRKBoDCdAFt6v5fXngPM3b2MuKgJsRcpZIsbuEa
I4901L50UNnF9iyM6+p5khaEdtQiALmUFM2S/VHN0cRQARRKzr82Bi3G2dLm4HRLK4+6VXQF30Zz
y98laLLLqa0EcljVRJQlXdQLheRKus2ndMDA9ilbJ0ACqjuCFY3BRDmv5MAkt2lBuw2WddpeBMn6
s3mlx4xi2kNGASPCZR05njDwpetlRQ9NrTgxewjUzD4uu5deWqVN4EZWLfqPlHCRGdYctdWe2qM3
MP5VYKM5BK49L5A6/nEV6DdA+A5LM/q50uQAS93f6NHLqdOe+im7MPjUkElOsBT7OU2nK+lw0MM5
jfj51SH4eZ3uH+BgoDMA8lG/5ek5XNvWaCJWKd3jfEedTGhhy7XEPWRb398osf9TDnk+ek95jVSP
j8rlzJCC7V4Gv0m+IKuaBtZsVoZ5jUb2nmWJIAa+H98uNLDPR+hdf6wZrxvH7ufoWCLrg6HqxF7f
M3quUckw04/653Ng69OcLniMeFcVLr4YQvxuHxgihmGriuYiyzoDCB7x3wL/uiDKzh21GOtd1DWw
BScIjl6wj4TEQ7Schon4v2prF/lmSvlSAgFex7TykErGiFoNGHa/PLlk9MStC8WCDBUYZgOhn3bD
Z/LTu0EknTVL3trXcY3oMvY6YYy/qr5kDk8fSrVs4zDiDbRgYw8uSMEaODcNGL7pYLqhhk/FfkCG
BGMeju9MHzZMUH+QoO/lwfjb0TaH4dEp2e+DVDcXcRFGY11sEZmtkmx/eZd4s3tGKz8p4U+QFxUd
RxV8WZeHrU0liKMut3zsSdfcLd7NTuAi9f8yeTj7r24uHs4fKpuZon0GJ+qVKNPidGzpxyl7j6hR
UDmrn3SZA37lPkv4xL50PHZFBFmL7x+DBQF8WO0ZEZTUTq3/hYOx1ecaUmsKCqSivXLX+J+/Cizq
kMnltrpeA2lGleClT9lQ/OKElJGUwNLJpMivX+nwIfdzd95I2mshmaHgVXKWBtyyLGqTiJXlcj9s
OzSfiVa/1tWT8GYoo2jUVbvlT4/ZMgoN9ciMi3VhQkSJBcqPOoLrzTHS7IhGoYl6tSl8xs+uRt2D
A+h6Fg+Ybf+mzaAkB2102Ync0i56qNJPWweZPJazwb/mHI/uPfAwp8BQVUkDnNjybytWmXWBmkOq
ISEldMPlBsbAes3dPr3T/c+8USI7hOoIEqvhbBw2es1WYKhyqlQlTq3TmU6WUqKWwB61e/uE8OCv
BHj5EF/e4+Vr5MUhXzgJoKVAwioCoxfoiyGH3tifyxBrS1PWv+DdlSF8DLfS0T6xd+asNklkR6Lk
Gy0uMTRAdzTk1X2cDBLQBN2AHSlyS4aUFpJg/WhsTwsjUxoVpGak//aOpDGmRPaTe+1ZXytPT74w
9PEHcymm90215T6f+qtrYvjh3+KRS/usr+ECJVR3c+J5r9/DqbpmG9PQGIL0+DU8ytPSAu3c82rI
3b1md4aUoeDQr4/nOb6Ctgrqtg+38QtCCLA1mbnoyiqlYkVCBryLr5jTjkBRuWiKzT2ty4UP0Qh9
HytTnvYMyg8J0GKEHw8+pAonWNFG9ShsSrLLZUHrTjfF2YOr1LHwwRQWycBGIBHaHWud2EjBQL+K
rpry+ThglWjenNI3OxtcI/G6Pa6OlCD4DMnnqbF1XgVIzoP0l7mUBYuSox69x2Ss+QThVDLZFTev
NZ5dKqUj8nt6j1ae0l4sSjnjQ4Ts03HlBXzJEne8BjluGfubR+PoXUNh5EN8NanTWJ0HAhWwVyYO
bYQZiyWrPke0p8bNNHUROJNehzT7s0ngAtomQzyIL5VW6ZJn9uaSYLrVdfKRU9Khj7L5WKfYzPAa
6I5Mw+4QG915SMsBwSgAaRHTQ0orxtWmd7MFqBHRc5H2fm8HIQPBpQvmeBDcjsJYe4NjO7eirXoy
7ITieAL2l8+pKZ9x6KID1SNTXGJSMlYzPXEpO2fkc7Z72MDaR4X9MozG2fqz4G+tU7YjjpFXMlrL
VTTYLPBr7m1SL0iqWKaMNtqf3LERrQ42DdIjY8EYZMj2Lf8fds3abdi+6Qfw6PfkBN+svtShPPIw
WYE8vj4YCSFmBvz2CdqP9N6PzKgdmlCsHzNt1h6QPbmlTcklHEVsR824fRZZmMbgmux4kcAJiQ7z
CKBOuc+gwn67mcBIkLqCxJkOfawxthGAXR2vhc/1t4NpRcdgh8GKQKWgyzPayTBDopXLF/EgCVy5
JNm72mB8iZDS2iDlveuRAZcQXgIGXUh3rIfSEIgPA6gOVUuhw5S1dtI/jr7A2wofkLvwJ0tfkMV4
aAKlaUzzZzEUrIGd/i8jTFbr7rmZlPk2pZ6JbcWmv+7DNGn1QikZNlgazkN8R8efWgNqMWsnYImw
md9AsMhfvV2toLQ3mNV/P4RLmeLz1jCXbWIPKCn26HcYbcceRDukH93c4Oaic1meRJtpxu2UGAEO
8j+DyAwwmnR9rdCs8GlqmROoHWBvDqzXYdB00rYrjiNCnnjrfwZF7+CuKaD6127QTXdjEWYrzSPj
X0qLtbEMmh8a85ttD1Is5K1u35ZDSvLf27jzH37mGa2/25ruWqH8lKlPV7N2SGJTMMBNauu/FrIP
JekQKahl97n8zRAw5jOkaZVK77or/xfEgwqDcTBuvbiHdQYMMmXllJqCf5ohpUa2/OGjNjTsmBwP
zS00W2lHMFpMp4LqLFpu6irozMo5QQYnrjTRi/vZrdOVGowTT13SFSNE//kQldfPEqbOZTa6UdnB
JnAJsByXz9OnIlLTIaGYynFUZqZjtTq47SomziXeTphFTkwjAt0+R9NJtWZErfIoj9aHdvk+GEuy
velVDgYg75clomB8cByEYVD5Lij9jTw51ahIA2sgwVwun+VtDfoQ/u52d5PnG9MJLgZd+UWffe6x
a4zuqGhNBjuJ2TuVrBvf7MmJVXf08pLox3nsF2AaqY+NHUVFiyKOGr4gB1GmTIdk9vd3tf3v459G
gXH84yRXuIs+8aiUjP0ButAaO4+Hok4t7QLs0+zfX3To8UaDHpHhvpDeLyz6XXqFFvv60Ra8VPGw
b+GdJptDLYF68BqPwmqz0cRHmyKxTLhb+Ko0T4zg6vw0oAlZjmrKG/25nvYB6W+1wf8PS4LOy8xS
BPDAItrj/c7LO/3atMBtopZXeOTPc/j5xtzYva91/27XOSK7arlZoNN3d8kujXaJOD/+0Yze6FQL
VxxJBmI2XeC5I/7SdxTOAdxMtDsudkmLH7SVatY2DPEy2vyTLr1RIKMqUCecvybqgmyT2e96NOtS
38tUrfdz3sWY47LfbrvJt2gUqgwL8rCLCrAya2nUwiSCka/oSUkwUfG2jMT9a4NiS3xChRXuMQ25
6sbnosZX5doaggonULazLRCY8IInGAvOUMlleoBnYuErNG7tFFv3rBOoezOnuEN47Trqa2iQ2k3z
pqujfHCU1Sz9bJi66UdugDoXmRJ28k+V3MQabd3BrPNASd5ugAOS+2KOyodfVDj7F639n6RyPdxZ
wUvU/FJIFdhDcQyRjZnUC9Mnyi5fGYSNnu09AjSCCeM8a+wStwxvvdqhl4CFy7/drRIMsNH1gaho
r40zHdebKXvlv3SvC5Moufppssmtv5Je5Y6VoI8tly/QoIsDJrZD3dJW2VeNG16DLNFRiGoGLM6j
ZRmeBnE+rj4oFatnR9VoUMzCMOMRQBIqrRbueCUVeDx6e3TRGZXZNf9tRBiOpMLlf0VUX6kUmiNT
oiwUrMhSsqnIBLkSfCj/mRzINF2vsJveJG/r39iQKRKxUIXdVhBtCcB8X5c6mhkAPO/Gi0Cx+rMm
MqUpyq7F+d1kgzLL8d28p3FdKtEsImC+/Kapkx7uut47GDe5GW4dvKk9Y3iIYAgf3rQLp9nDq4Ma
WQ3W4z0GAABrMVX8EV/VAc7Ap7wS5DalJfr1eMpK8ZtCEJ07Xx9BDV2C9YUpPhgJ/iJSFSqjRhXY
eErvz0kthGKm4MG5H/BsFIHVpR0HsAwrZklNo6Hto6csqXahberSxXTbuPKuyqU3NAmCFvgVITaV
tskRyyZYHLmdJSyywhpHQAm6I0nQJWB+3NA9AU/TZXdTdR1aOMOCG0PhDYxU83GISKXifKBfZBWT
hLV+Bj3b80TLNNnYPDFMXCq1rxiTTQghWrBzZ04KggwqorB9CqOKV+baxm8fDAcUwvST0zeAwQ4L
G7kH848Gsstw/IzYfkSJ0LzF+lkkRD6w/l0Esl+jXmHwetGBZrnFVlW19HXydkYjmqPgJn+QFe24
CuMTX7p9cHHDMvH9+S38x3s7ifA2kobuUEkz6OH7QVy5Lqa1zo/XpK1nG7N8tAO/cPAOJuVLr6j4
D3pMdN6qPzwKT7E7DeySrFpn3IodxN/e7yKZfwjGxNNH+vbkQLAjpy8d/crsn512xSwVuJhCCcoL
oejnSuy8WYgu6HjWUUvsrhYG7564UjiWZXGp6cwTGTxJMpvqWV2Bx4zPtT6MI1xarpqHCy7cSQ6H
f/pNJg5PWCG/HM/Z5T984dgBP8jkM5DoEj9eUgn2d29MgsmUw6YlwOfDZxpPjWZMFjOvgGObx6WG
JwJezgWLo0Wih/w9AmN2by0phYPAdiuHyjeqLBH2YdJ3bTpvE2rpUsq4c3mTQVXPetB2bNxK3bLB
5apBUaqK+YVPgC5mdOH8v8j8bjqxPPTozLQAUmQynq+FkGBY6pRYQ5z+7de5LSGZ3L9scRGphwOo
nHU5uc+p0/6XByRw6H9kUL3xTGr89uQtvpj7hlKiWX7JOK1WzJGBD7lbli9FCSIM5quDAM6zXZKX
NZ0SbLZbPUJBfRvKl26hKUZix5DmkDHiI+hegczBdfsyVBDUkNlQPnercdIMJs8wjuApmFTfuyO3
EUUtcFYIM6x7M8ZkYQyLgnxIKaEBBQoyS7SoCAGENDRoMqJrdq0BYivTscCbTjh3XiEhXxQeNHfR
vPusfLFA9HUB5Ou6M4JHhP6pCbkZ0m7Or+oHFzQnUALHOKhRvXRCRU/oVgUkFhgUP+OXjSeYY04Y
qsgTCW+/3cJzJWUfrNiRqpnJgjIAwTSITyVkDMbbT7molSvzzk0773tdGgS4a975rYDp4z1FQT/g
x+1+t349fyh5E1sBYLDbzwV7oTeDQzal6uLMrV18O0/UJ/VCBcGrRi/sFveIYJ3Nttn26BQRQXTd
iRUDHq7jeJijdUGtYmvMur1BtJw0gKJG9RoRb3HOCR5Tq0mxp7XmxHRB58I9ZOaPYyxAXam/ea1E
hH1GXvnhT31XFxMzdTi98AmeUcf1um3zqXerYNIAlbA/V4/WuNANmdoVOoWv0iKuEeOElOUnJHWR
jguYW4RYPQOpC2yHgTwxGZC15NoKGcJ4S+DddCzLjByrA9X7JN6KS/O3ZN4WMEH1TjX2VhilAZ2F
vywaOJyZAop+KIKSQmXlq4iC/vWgtlH1UrW67LaET5ofoE2Ue5ErxUuqMOFaTfQ9NlTx+jnc9/iq
GEdGS8A81fNWw+/Q1EjPK9+0y9c+FJpumlLPHAd1btuicWGxTnU6QVNGsDbaAg+ubupI4GWCi1at
9eM96GPMdhbJYIbHDyvojK2hkCA3E0mvKFrP402DHsk/QubzhrR5R8ghogu+jplZ4FWIwNr1/JuT
na7SQWlO1tgBs1Tr77IT3R0xNo56yM3rOC7+sA+c7KquirmtfgUsYNgRTLaPzUCbXwHTC9eQLfuM
hUUTeWNykcSI9mseYWDksbShRQAPLP4oNlsiIE88eb1xj9Rpq27F+hQUacAvZCSYrF+eQlToze63
5EMmEt1ZT3at/MiUsnslyfzJB07O2rut+/jyi9l1lW4TuesvS+OZh5RhdOizaIQMjxGMuGXgzSbG
lkr+WBeJXJleyRvR4KbFztHXDJF9SAiDGCQYkQtbi3+ZMW+GNLu1rvtDbpB1pnsHSRAGDeQB4dei
rD/YyyiqViuWUoq33CZRxK6owMqrVYcvKSwoBMkcfnWoNOdgzPjNThWd4fbBwADAp5tju5+KIfaD
FBnU+z4WShar7P412Qrh3BjNUKlgHcVzInis/rKRMBsiCISto9+patvtWFld27qj/f5NPLVNkRTl
xqpqYNysF911CYiA9vnj6tfepOKJU0Pb3I7DybJaGBRKAPo4Gq/jP6Xd7vRPUv8J264dUzG6/+kk
71F40cMT61RGkA2wTNcQPcHAW+uc5BWqo8i/YyP6VFrob7FOloLs2DnlMo7mJ35TC00GZqUCxro5
GusM1iRtfdqb3wJajdkbDulCeYtC3qzo1Nn36sG7UUpiAV7ky2GqsZpAAlT1qc1+fSpmD2114GVy
nhoKQx6pK1+b8WHdowyjHaRAPyS9oSDYP4OVUC30/cqnAhTY/N0mAuHbpa5kHKGm0ss21vhZHGrH
DivNoeoKtsYR7RVOyIwPWTVI7FFYvC0EwkVuSjd12dwyyV3ustFdDMYNcFY16QtVGK5PzaTmcAVc
95U8uBGR3G+AmuCHbe4O+UUUcCsFDPPCPllZqY5G0Kx/3ex+Udi21cEOqY4pYEIyRIXJ2kuHq1iC
rXRQdXPydJ1Z6uIz+SOeKD+DpSuzpdjRCjkmhPXukZLg2P4TQhhoTuofN7dq35OS1nLVqS3+cnHy
ZP9/69Yj43+Zs7DeKW4s8itaikzFeE/J5GuVLKCyqqOVps2KwSaLAYFSmkOT3bRwsC8QzRLYR8G+
9BDg6MAb/L+UJugXPQoSPQVHW3HZKSmtgZP19mWeLTsU5oJ4aoqG9Xy4p5+6yrRJxO5yNvlHO5yl
l98ktcM9dTjiD9vFsE5PBbFtTO0vzwB7nC7q+Z0pUZorNMWlUhp8hJ8H3jPKo3/BLzArrGB/MvNH
1pZ+n4Ia+wB7lc4pFsN+Ve3+SNout37T/p9SEIw8eGKhwrcljp39a76d8QBwCBhqOmFppNRckULe
IoNmiRQA2ruIyPSJIQl/DWGp4W1UmXiXOABvcACbuDUjFqi8TQ6MuqDT80s1j9ZQGLTXroYvUXUY
k/XJ6b3YSWVMOclfbRyH05/flZzVeELh8zh1B+p8s4hySG58wxumzl9p2X9l5+4SUi1c13X1yUwc
hwHcE0ih3AMmdCrhd0U5tqDCuZimcJIsq/QJplAAHF26/6+vF4JI43i7WrqSGTx06KburDH5IxYs
l9NpEDNIk+lCLUbPSanHJDDj7/AfTkQCjuUkGtKw3nTj0Ji/jReUoGkZWiIYQwQ6X7sUHpc48FcM
dfbX/v9z/MzLH6+S5YQHdps7TlXS/qpXGrogLSp446hy/z55SD/AtXWcsEjctmeyO0AAM8BAaQkz
q1Hs8o26pNbG/dOr7uWTsOdm3Q4tbOBIu/NKRQLyRLTufVrjSDWZ0HFixOzmJrxsGmL9BGDx2jiy
ZfdyKNdq0dlZG9B6zzY4G+hHGGb1j835xOdK+FDXxZzckx76SC5k6Yplb9GI4A4cZVvkn62I4m3P
c+dl1Mxdz3+ROvzilFAgSBHStAVomzs0s1+y3tkgVnB/ltGVaYY8zTIM6yQWngNM4VJM24Drr3Zc
xAtPb3JB587gNAFAEynp6aGWabo12ZE04zVA5PrtkqLyqufYhyJSOdP6eRhLsqifbj3ek4FMyhaN
eCW0t1RMJU3sCDz/T3I1sH4ySKzCUCC+v4aDzcoG3rRNlym8x8fY+HaI03WG1y0kWSTmXyo91wgU
I+6aJL8h9FZAYGX8Hf8zSL2fAHWto0fXad3hFRcJKG2RQicc68kqItotQ95cJz+gyg0M7tHxqKaX
NiBdEU18o9IzYzXI0Gmq4pr2/q5y1fe1+Leu4ZWV5msdwIWAV39Bj8Of3QoHenE+bG6L/xvv6WHV
lMKjQKd0it581Uj6Mm0Un5CxvrrWdsQdvxCKvFBc8A77K0avh3YmRAWxASpXShQ9I0uaUAR+CVl2
ZJ/RnJjDF8yNpMWWm3hH/UuXupNcyTZoW219l6/sB/Af98aBdBErQ0jneBE90SsDyhWSURrge6FI
UmsvJdMFyHDV6gHaeFQBvJfj6WFnlygAQt1eT6np9vH4gXymE8Mu5I17VioQpif/lXGGGnPyrwV1
UZFNjnAiK0L4KSf7LNRlRNSuk1K8lpQGdsfJOuKzD+4puVMWJEfw6ZZom4ZQm+fo3/Pua4+7uULv
aiLIVB4+7J+MxLV7ZttNfasbP5xTx7rGN7LsDrMsEzOpaYkrkxcXc8igCy2y7zKPQAi0BNX88pgw
EqbT1Lmp75KjIYVt7UJwpJ0JyE1VR2IS/isCLDw8SbeMqJ+TRgYzriIb08/j+bGjxbffphikVxyP
IQOUAK10lfJhr2Wzmn1EaoBgXUO4JF0twJ43+9yGpWVs9qNTxEpMt8hH5OF54qtiWfY4Bj9DQiLM
Bi8C0GI83qr2ISPcvnAliOFsUgEiRzx2VXKJyxbJgdWIwx9DchKngMlSThqm1AJrREdObwNILYtK
fYv5j7tRDTLgUsDYZdDFLOIevlfAXy7Q8Caa4NOi6uFeplxUx7w0N0/bJhW8nQTlwGIba2awjfid
VybPgo8LuO1Ur+3X5pzXw266B4fpvVj7hxnalUn3uUAh0m0pmUAkbmZNLNLkxiwg3NmteHDBNXX/
Zvx7FFhfHedI/GxyhTfvpleqDjkSTUE+djzgHR3BAGPgWGTdZ2Z0t2VInMqNv0vhNWKDXlOi27DI
GWCzC8mtFfBQ7RZIR458phhmlIJF3wawDqtWuKbU2TTVNBNkqSEZ52677H58C5fzkvqY5lCrVV67
7/qBYeZZbH5dtLf0FmhTF4sbUlkRgeNHGcfZ/zloaY0HEwRza2h5yz5AMSGw/Q2DBrzJMmRlul8C
YjftJsf3dnxvwtL8THEavB5peS+MenLEwtP62pVqIqXngSuNWfMKOT7okDqnvQ+kJ+QlGO1miTov
szEvTb+ZtmiDJzsfK8mZpHyD27pyBWuKE0xfOfhbUPZVR+oGwSMrFJqSmH7PRn/C+i0L9Yc8VwWE
yOJ+2pK04a6qpYbhMcZfGzzfSp3D0ad7Xh0tZKNftEVe01R7p9xvqXPn5TjxyMhheHfgfRLQqgWG
OS+e3fRCwrBnOvP5YXBcPlN1Qv/X905FIEA69Ssyj8/A+RawK/E5YgmLMxCYagbSkr2xsRkw2skF
Swtxn1Hcexln9JSGd69SSnwBtMMsZ1xltOEUUObZH4o6pqIBUetwvaxX6azirugKLPErpLGWWxMg
hW6E7DZV0VB69H+vxurjwO3LYjTaH34PQfnigmde/Ch2gKsAWPc9bKhoorOEZ7y2dnQH2F2E0WoI
ZDW/LDAjvFCT9QkSm+86mc+6hBtA4xwIYwXokDNpAb0WQhaB5GlSk26stvMjmnIwMUuryjrVRFYw
WFqTJ2icTigQ65dJcTG4bzktFocEESZkWn/aQZvHKEJ0by1GrELsNKJo9iAPNnJ/Fo1k0Wvf4noY
AuhElooMVVICHurbOoA9E6234UROCW2w8LPYCc1pmkAcLy11p2A1ZM8YR1y8t0lCGtNApm+nUcyP
f2m0Nxpo4V2qAYQ2mJcexZKAOibFRMRh9w3nPVb0mWJukeN3MQaeRpHpKkcZRtzPw3hOdQkbpSDg
RTkt6aTIkcNizkkxKCRcqpQjlCoSQMT886uRLS+Ns6ITjn2yC7Hv0NnFnzW3SzaTCeniY2TnVnNh
xePNC2rTonOIyEMaw+DZrBULadteCu+sAw/9fChswM/YjuCGerMjb5aTzeeyrR49MB0pOBu06iSI
LatDgQeqoLiklZL6FzQZ1RlSqIChYml/EJcrhEFXHsi9vRLsV+K6sDqnGsBKh/vYBJAhaHYFDFcs
S8jrFJ9BERoGbZW4473JIR0cBxbi/XQRMTS3eqzBiIafohXcqAJsc0ZKMP/sgBaO5t939VSIXG8a
unsjpm4LE2dnijkfCaLQ36Fyp5i5vHsNsC6+2TkoCeaKLqjWgT1TaJHD6ssfcMYZqBH3UcTy3ZjH
tgMXUbllKsWeLs0vEldHUOqa82DGDbbuZFOmHxHHwk5CQ6cZ9ZFBEx8ZVslL+FUkUJ9twwmaZ/vG
yzqzJpsrvNT+4sCL4rAzxuRVquOuvUExhScDlJErxsL/zg4LcZej8oCfSuwkHJHjb5wRkpHGnEjv
jsCoGhgeyWn1h/evUoR0YgvQQoCUzUGzEdzGb4Kj8RHcd1Pa8gjsBRn/BB2T1nbGVb5s9OtW2Aow
ApnxnL3Uy6VPKIhIjxxZF+BEMQAxFayCx+8qfNGP/Paxhf/MCYIq44M884zZ7huudVgNNE4YY59S
e17aPvneT4K0yXEyHzZNYWCJX5uluXb2l8GLwj0uEBRcMDcUoobx6XZuan1y+iYNhRkU3FmnOb2L
hhUp/o5bVvj5tDcs6tF6lhheXgdkq5WVKvrVaStCDnI2o0j1icjbSoCWS/hpByDtJxhtaJKWRLua
bOCs3DoDe3q0q6vYYuRqQnDE26jr5LW5m1y0Cy7SN8ZznOvyIQGJmUZYtrGl1r8zzZk3KCe1w52j
NOK5P7m9TfLQmBcfJEwdaRo5NQ9VOIUSWOipmZCjOnp/AvqWlscInAKSsDbtru4n8JrUz9d8uQfH
Z/qjALniWoYHrgaAj3Nx7J257efurbpSo3JOxPl/CvvP3DOgYtXCGZNOTgqu1AWrlgFDrSCYN8Rg
/s0IIWfZqvvTy87tjI1Kcbiea9YigaEpul4Y/ysdnqqP2vMmhnfnISKJ0lP0McTOa58KbaZlkQ/4
4ikrBrOmqveW+zy8qHv6YzgtN23tpKUNBy7ef4ELXt97p6LDwr+6WzibZ4PS7y3wRtDeXS4V57rJ
mU/y7ImssLGvse8pSC8RWpQTzzJkVbd5FqWKQM9wdXRjsUFmmzkhZaMTPyQC1cayhHGX/vRmqWiK
xhhDb5RYXr2I2Y8AOgrf+dnTCX8Hdj+7XxY0o7Jn3iSgNdLsgUA2AGIwqSIcDklediQd/GPoQPBx
CNTda16ntVmDcLxRPiPCbtMdgv9OEISERPDHMZs1DJISyZIGrmqPLoqSj0m1807mJtQUoa0V+AQH
qtBgyDT5CE01RutrYFIbL+0296MH7/GMOb+Q5v+uVHOV5psGQzJlW2peZWTnkJtWFueHLUYxTs98
/sbnCqykopcaHu4d8mFL7S7WbvVwUhl9TFbbxh5E+qdzBumpg7YMxdeMc97zfLauFIaOgGOr8D15
50bAzeePpAdf211ac+IL/k2h/OdsocJGseg8ONJFYRMcW+KmWwtRuLXc0jgkpz2gEqtYlxvOYTCQ
i9YntS8NOlB7cgSg4BXUnO6lfDQMbF0F5KaIytxllPGX4IZuQKOxwzTnfe70HpF6tSOFXX2NPsC+
tdFddIKieDb9hSjTEf8oG9YqOp/IZ+HWhVFc65VrbhBcDCj5ladJvI8wzAef9jdoxDPQ8beJ5rlB
eByNlgjIc82L6sFmfYKb2EuolGI1WDJMZmmihGwL7aGoVZRQM7MufERFG4kaD4zVmzgMetmjlVVk
6GyMKQlm5enhvUgNQP9R00+22UG/xMAJg8ICndwsD/HeeeQjbRc6FLVWzKc6LZYE0L0LpHFySWAQ
qLg0fDkmlAO6ImGZjROj3kZ4XKeUgmOd51jZ4s7fmoSs/QR5ASqTIhFzvOzB9KndJJXVFQWL4rdI
znnSDDCsCLB/pDCjv4BGWwD+Ry/3PUZ0wj0IViEoovloHWalkNt/ctBHKfeNKDXvJDvDq4P9px5/
YwAXAUc2XWdiIc3ctb845qL42ui5H6qpHk6p75JLVI5DQHFmbDI9J+bCYU747JeNxL+vZzHsLpsx
5XeDRGU65u9KkOvQ6pCFoa79FlwpYZIXe7A+qi8RYWTEz9A05HmlFUakfvLcmL+ANKGdjJ11YGV1
kwq4mPbz0qVSNACbajsB5DXiPxORaTSHOvOYF8pW0QEfuUS6ucfuHKBEfiXb21eziZ2zjdVo4ahi
/Idw1s0HFOve7f4w3ENDUrLoo+xDhHBnWcfplmB0kz6JJTIpDz69ED7wQee7KQC476qj2igJxrzG
l7mN++BaKNA/ZYl4aCItuRMkFLsbiIizIA+6IHYjgwg7gXgIP4WxdcqNwkjlls6rbzWa+exP+WpV
17nDv6ab1D1tGxtZ74AlNb29D8Ikc/CMWkfJrBwfruEx/QnU83hokF2zXzxdEBf0U6O/oY43nygU
yFJAwdQErHXeIX+AdvsEF9ER2S+c0oXIpJovAeDlqn/39O4N1scTBnqpFSCH7DgkXMOq8WV6Qih7
kRYCFDGJlDPNqtxNr3+o6yrGYAX5ydEnLz55UsjvNLEaNAwIQgo3VGV2HtBSbaOWasl5CPoSDVyF
RLSoYogN1KE5MGzNUIjieUmHYcBWl+VQ8Wi9Lm+4WLpYgJkZK7Rg1WiUh5QLe+CIs7BcFXIdxQUi
z92o+nKP6mQlRrzi/nKSJyddjitkpZwTWkdLsZ3/f7j3Aw/1ocIpxbAkRV3W1H592l0jeAxWe+eW
fuC3imAVlAixOj/jRbK/6lU2D71ZDizIJjE2mvm1IW8OVIqxD4J4VIBBNw0igJ+ccZUftbrpiLkJ
mHAT8oHIXU8YtmoT7ElFlO0efAsSX/lDbsw1/KnFUaT6ahjBgUtCjDWI1g8QWGmzJMFBSawMZNBC
hULTHkCuYHXETvKgE0xFLSv91w6TtCV7JKGYN0MfNCGNRJwrHyHDzU+sU7jmjbneMug2uh/As2MM
pc57FKLLn1Gp4ZJ1msdC/LSSyTKwkGiIdDG+Up4YG0NISi3ueJChF6Czwj40qUcVEnBDrtnM9eY8
ohVXGy89CyphUkeEcVH9fESBQ0Poryv/3skyKM4UW5uD19x16v3ZNilrTcWflB5159Mjy+H/A6y6
sy+Q+NkIwgsy1V1fOYDAGMGxBy3Is/s8V3seqMmfTLsG4wq7Y9OukDZ1E9tk0UOXllYo4tB3Z/QD
iZllEGW38++ssIkxvIxC7wtB04m2c/79kwC6qSUVKziwRQtMk4hMrL7e1vGzgo9xTJv0iBUbxdEy
JG68wm/6+ELQBY4n8VkWyGeEetS1i9sdWeOBg7UNAYG5Y++pU3IP9r19rlkLBkLM68Xk7LuzfQEC
1Zyp+NKoWagX8ul1Q9XFZ/u6/wiDQlGAlTYsPwIsstpd5oXHYjhVHlCVD21xND65y18iR61JUGf3
4JQbkZ8mffQ+I/BmqCLxNNZ3KYoWbGNr2SH45V6dY7/lJSNmchKLb3L7UlWS+6IgaeC6irz34lXZ
pfJ2eSFlbJD1s1RTWRgXpmLEUFUDpV0EDt4JB9HJLFKVWS1kgfyDwnuOLHJ0sCXh7+DKxfbKgizu
MIAYkjjqU4OsMOUopk25jFsHg5PZr0IuPe4ekV4M3z6vp6x8Xgb93r0Bt9C4xU4By7AoUAyweAAh
7H4ENcn7vTyzm9PKDwgRpApGu6xcbsgHUmw8Zn+URyam63fULXTWGB0zIhHeqPfYdZ9RbeW3EpX9
oOhYKlGaVAA2aeQ0iThQW2ySxT+1eQE53zNzTrg0Sxga2LkLZKC74j4dKkWzA058/FYqywSRnxmJ
eaabkm2sYIBPjwV9EiAdYEU2qnt3jYJSSWZLg3xvik1vBbQDFdytMm8zpXLwwGlfUl/YVlREeLC7
oImS8SX138fwe76VSB9ZQfk/yWK0fEBJ/uugQLDXB8WwuQ3mwTQqykEkeBN1hXEcExZfU7JbgCxK
2sM3iU9dWbTIiWAhLW7KEaZgr0wX56cVJDL6y2o8xZYweuaHxnmiLCUahF2Lo/au7nXospO0hbV3
4CH2vkM+jyQSresg5Qezn8NXrpNA5ZwlbCm2emLP/hZbKPx3Qm2ZpOoke8CnGXvOytmdlCDpOC5x
+mYMvjnA/K6HZz8Iy24sToVAaoxFlDdG/NHKZ9g1xAszOsk9hNyyPYXDmcsSEQOVGBlqQCd2lbtH
FBIapCB4UDBvwHNGP20NoK4f2MZy6YsGKGQaxqKvlaqHQDZ3qFMp5y5RB9r7oh8jd8mstVrw3VbP
C3iH264wS8t98kdzwB+9ai8Sk0fZZ0qG9UieJf7+H/k76YMuXpm8/pFk6I1ayDLovcPGjuOBWEaA
aJ6NVRiXzNl8wlkerIJ5MHrVbxu2S4sJypNdCTwSUZefo51tV346ZzhmqOu5Xs08lKQHhuwAffIa
wZ7bG3NLL65eu0pJ9r3461ij8s1gCJO0s+UHAHLYuCSfWMWgR26drhqhO7M4YGW3Dgaof4SKB4Zp
fendqKRKUsrC1uRHoLETRAe9iorlC1B2qmRs0TvGf/Qn9qHcnNqM5vqq+52LnOFaRF7vVanIHmVz
lGmdO4NJQ7mJj74qBAlkuCL91ZvX58ORT810nkTto4+IAsyU+9RYvkl4v5hrkKzJu4M4xha12OTy
MEPSFnQXNxOjJvkJ8VzjVaGkoWlcqQ6ysRWOGJLlgFfnigaPX93m4pcBAJL+LY+0ZVo9UrPM9yCX
6LQDhSNa0WgDGMtcKyKkZ2HoVBT3VqHEWrqRG4qR4xj9FMGENKFbT3qrakneLgEb1hm4tWhBkmP0
h2C10OOfWA74RXLox1dwTUG2BBBQz2rhgGeY2ma1Bcq+TDdUOpLYabdsSXvgRTAOdSK8sNTlubGf
zHVmVtLLg9akJOH+tP5HBWGN4sfZAQSOzVsBTf9n1943WB17Dj3rPYeNQ3juY6vfSA/jtFmSbfIC
4iPCUxzjn48GTkjUF28jjHTrqaqBCtEuqTJR+7y7PxFhlknxMX1KEj0aX7WOiDC/ynfb9jCz3b3Q
6Ibvh6zg3kgpz5oPQwBePSnRlhWlz/3indV9upt6RlQYoAzSiiDqkqLiIyeLUZWaKcc0DxcYdI7z
ajUVvvUTzOJCdpxqGNQblC3zMUF3uBh27Wj+Z5KHuimOBAns5EEomZH3U3mpfq/inMMxW+ToDiJf
rLz4FzqxMJKNCuBKofnBbr86CCzIdjQWhrzJl+tFpysbcyqHLiSk2RVHra5tV+qtgvdi7IKnW5+O
X1IRtwjigk++Od8u8n9g3rI4iZ2PEytHNGjXC6cuUUtE8fAJiok7cy1e/0p1vuMNQeQVyyOe4102
d5WHiZDKUP5jAQV6wli7xYUcgYMO+KKboQpDdInlUm3/Y0zKRr/zM5s7KxSvrfPPuvZqmIpqJy6g
DchFh9B6Cgx47OaAPbPugKU7zNynQ/pA7Ekl2VSjywKCAUcn5c7/RjkanShgCHy4jhgfk9Wm4VcP
lb+4xwHINuUnyKluPifX3y8yW+Gv2OoW0aQFL+Ld/GaATwDcim8DG64kJdj8u1vl956pL9O+bj0e
kNnGIJxS38qwzxnnww0JzVcZCaKfIQhX/aMJrLJweTw5pK9qbU6XN9CL2ikVJZ5oeSGe+h8Rtf2D
UgJ9hAe88lpTcLP20iq8NCtwVwtX61ZL/GHfK5RI04lKDPFNN63sSXp6W8RdqZ4ck16gg4laTKMl
ysfRAmDq1+jnrdh8qgMebNmqHJyIR1Nue62aXn/mM5Rv1JjYw/1FbuxYpLuy1jJnPeo3PIbUGaKf
Dgmk5y5D+sdiw+1FjNrgS19XkPulwHKbilFHkn18RQIHdMGZRk/nOLQLiJF2QY/DOvoHHqHdC7kA
BnMJ7rwB2gi2ZAeGf00vj7GHyGLwJRSrZEAGgTb1/H+vjjug0HCTzUszU51DngmM5BNJG59oUH9I
klEVF2CY1fgMarl/sgxZVIGWtnthGMh+5x7Bs7OfVR5SSoZg1rDdlRskvznNo+kewvAbtWMkZMCY
bZq3i8Q8I+2U+iLlZHhgxItQMdtZJPskwzZROVHE1hl3nA2lSLNxX6/jHVI4BqM8/ki2sh1t5Vyj
+ffJYeo600V4uHcwf9zl46M+qBEZMPoH62V5mg+epA75ot6VmKnajIImt532LaSqMHqLq9utdveQ
fXIpuhDwJrMH6R/mthd9W2bpLoS7JrMI10CrGSMSr/vJwAz3o6Ia6qleoIm4Ib1UOUje/RaAidTE
2I3S4r3hoGR03FOppacPNNBBYFlot1VneHJiYShPBAatyte9omtI6Y4CA+C38eI8LrKnXvJRZmuO
QYQmbNiBU8igBkbrtDMjdY+ldxcWduVZBmQKo/J+LKxoO4UEe1QWNEQsSBpf2iy+wxHs/Ii/kHVw
PvDDaSDohc6yTH2bNKDE0iNkn9psRprduTBVh6uQSfA3gWAQeEyzT9uFCvMdlkL6RNVcf2zxxpJC
Fcd5NnULQI23q+QyHZKZQBiiBQMwhanGNUarwu4NnctFGljmpI6wNptgcmQrSp3zf3clbWrjSnrN
T5P59VoKAZ0d49iRkQKvdoMhk86ei2V8VOqexKXKE3QieO1t1LJ0WNodVlTRcJcWuYp8Ugqex5U/
Kvb/+EoCd8Pe1M4i8vLGnhXWLf5Q6rmzQ/GYQMCg5Psd4rFTLAXbid6kxyh6Bf47Xedn558N9yKb
FqggFiSn6v1PWu/w0wVMzxRWHjTWH4toRxlFOk0jc/p4ZmPebaO0jKSlvEp2IbBfYPuBhG6FK7bv
m6oAgkNW1PlilEShSIA1Y1odda0txSoaZXkm8Rrer0CxR3PrGbSWS7Bv/cmGf1ebPiXOVXUpo/o1
JrXGlztDYU1lGIX2CS7P18TuquybPgJMlXl7eI4kLROaPb7HanJyT39xoBTGW2roYiHxT58frUD4
Nxpmdb6ucmxciAlaTsHe+gyvSXHjYLz4B1hTdLUAcz9KCYAGQpfleL8JuSkwmxCNQbiLv8KVx2GY
EtmHrjAwD8Uw9PoxL8YjwNyZr5fnob0VbQBpNEVkhi84APi2Y1xoBcXPcoCkgq6dIR1VgfpxS+Su
TMGdpgBSfvusfhhccXrGTMZBkZM7S2WeMWiuCkg0aOqUj6lNXgllyE0EfLxXbWTPhq/bzuAKXpz0
DrG1V965zZfwNlHhuITArPFcGWQQxPRZuhadv3C5Pxmu0UI9nSFOMqa3vCEjLjBpTAA3lb9qN/zl
AUigb5jAuxyRu14Nf78OTnVavr2DndyLaN5aACBYZozdk08dN/q6ARVkn8jHWKvI1IlepTwkMxOA
WyGO7Mc/TZf8IdipqhGAN7gNatzxZfe701IMSCqr2ls960I4etN5R/MsDFOX4YVoVT2/X+8Yqgml
jYUsn/wzwntHATJcdVt9/AVknL9+dCtYJ1YjdNHw/uJ7UAVvMhVo6cD3cGWtayQOjq9BucrV/430
K5r+qpiOKHf4YpvVjOzVGApUfjBCJz+5kq/GrYpA8Z3mvNW1A9UI3dDPOXN6ahPmyin32XR8Fdau
3wOTYEFu3ib8wKefyPLTvlHHE5kDnDNFzkDise30EeO1RmCsVfPZu2hufxrVcKLcQdjAw7stCy6y
ljApCa5v06ph+vNslxK1C6dDcEfQBTpbBuhVkdvkduPXKv85gqR7tjQNlEOIHIFu5IocAJPt6mkZ
bJzfyYz4b2NV6ksrowK9immKnobeqBfue/Sw7XNvxwqkD0CpGC8qeLzrmxscSTt8aOJqpfhdgS8x
oIgkCVuL94XeW7EfTSjo/stQ/bop2NG0nBy1k78iDeEwirtkPkoLFM85bxR16EIhMOPG4Sgp3MDi
5+XM+Juh4f4JOrKFhRtH7dthYdaqbvl0bzwr8INhqmXpGHvFXsgZG1jHhCwD60vprKHRsuOsUhtZ
f5H3mgPh8h2ybXMDfc9iNjApi4w7inFJV0skOThfFLpUQDJVntzz1Bt5y6d6yGPWNXfNFJlVS7G/
AQ2dkcZttFNlN3gijd7won8NoMiiLHos55OY+k2oDrUTyDzh1o8VWXW65AbXi8P8plPnVjhGHhCB
vWEGtjbtlPwnxlhAE/2lkMyrG4lqh1qXlR5egGQPyQ0cwsbneU9bquWJ8IBX3z6jMf4fa4X8IHSX
74VXHdpZmQlEtsU39mehP90ru1HNaaFNhrszm4Oifejsub9+yzlntkDX9Fxu9LiJ306nEz8iFdhn
Y0wV9bAzquNMy9ojdRQhy9Ob0iy+8mWm2hniSDJfpRf0NHgtS+wmWf3zncJaA/Agpr7tKgQxtzLa
5+bPhO3GO8yE47lhpagu4lkTwIqF5/0DPw6BgA17mUgweLLzw8L6SPRpHG2klHM6AfUivcowPPWO
kWl1BrT/Dw9+XxL20Uv92dgBNO39w6XOBcqFlY1senG0POjshzUSWsGzw21GuYDvbJI7SrGI9icc
R6L+JRVrPS9AN9c1gJqzz3Wo38A0tVCUzPVdymt4nSt6My/99XZZpuSRh/7fvxg56a7pA5I1D6No
UXTIMTHC97jemmMNRPpenZzUd8AaFc5TT7Hl+wXqpMepxE/g2GioZJpD597Wuz61f1mjC30MpNH5
JDLtOewqomqJrfroPtca1y/eXaZEqbzJQ0+9V3ITh6wTerqG/W22QgquaeLusrmcj+1U9kDDlqpZ
r2yHS+i6qLQlAvB5thD8h/YBk8WjLin5Jihupl/XH+FFxQWUZSG0y8AkNPMytxw0fra3nPNjD+Ld
mUfLVm3uki8cvLx9WumEhuHqUguEuLT0PeCMpXKj5rvDKTjt+aFP7x+aI3gldQ+GGS8ycLhPc5VB
bsVXVAPyiA0BmK8PZ0lVMzueB7eWXIrSd9ba3QMwO02EVablvtuJURlk3BTAfiVRMuI68iPjFTRl
hq5XjNog/VYjoZ4dgMgYSSRMXKOh/cXoDUp8gH/kMAO+3zPYwOCCDgkCglNtgtgz7lCKDlvMt24x
gS/+r/bCiWoN+FCLjlQKi8llKn3XyI1d3elgETIMmZe489+1dbon2pLzUhb9U8yuiE67uzinAqcG
s8g1d8yisqwMVOHcBeOR3bXybY6RnkjaZerPK61LvK+MHTFf12k5iyNPYm3qLl0n7ypaxqmtlR6w
xoXJty7tKt9pOX4bidwYkUZY2FASoqneujCVIkcSab7UCgulrjJDYTiIXiqhtc2z3cRTV1oLMMU7
frYaYP1taiYquyMwiT+62AXIkcj5GIUm1AHCV76uLoKvwMQHBRaoM2OhD0cdPIxVEexIel7tnCEN
edVNKzXpAfCtM0cygsHDWp3I+1V61hCUQdUguCpZKoFXhh2Ihni5TT89HNMn2XS6Mo1CvcQASS6Q
hvzUlItqBPoU3nyPQm2CMEa5VDvKRCJfcTCdqTwEMFYKoRIlFWIhSx0xMRp8GEgs7vmMbck2goMF
MmCRpMTwJ/zalk5mykf1Os+uDKmsL1HXnzFSkzNPlBqMCyP+U75DveNEpFJEJymRvNsbQg5G1xoZ
ZhmtoPFyK4g/Fjdcqp72uhQDWrPJJU+si0BQ2poGq/0PZNTDbQmiL5kkYVdpbOHg5LdyOxpA1sEq
bw6oKHLe/y1msaFSyJ673SgxyaM/soNzeopoe+X8cdWlIp7b7hU/UVf3oDStP90CEC4gTWVuYbzV
x+5GQTq5Dp75uxLEDK2es9tSSGIyWA3QlWQQnx+fROCtbHs+i0bVzVuPjp2vMBvnh/okE2PHxing
11GAG4vrqkthLy8q+d/TAZaJ1yoHMVUjxffnZ4b0KsOCs0jZs6++nf2YV7bTHlb0M7XzCcBxv4Yu
RP19+NC5EXScQ4uUBZJ5TAJcFIpJIHilJU9N9jIigEVT6NYC+jLnUrmV6b2M6MpFyKzMcr9I42I7
72uNFWwk7oov/pgx056/2CtjdaatNoFoKgPu+rFonZ0Vk0Pml7hKcVE8RMBuw7cPU4pVFdUIDT9I
koBl7Cy2kqVdIFiJSI6xHvxyFUw+zAgW1Po42nSEdyepsQ7710ssIkO4yhP6TpaSuT1OSIfL92ot
ygJMmSiXhYPZFuy+YLc5hMiAtN3DRyebgURjlNaR0A9oX/SehoQFfbELEC4NGsqxST048LjqO0Fw
uqBABG+lqOIh7S2/rjKxY8RaGTTYcGQyOiJUa2w8BCt9DZM1L/pwgBTD+Ht/t7IDtWanRhaXHb8J
rdquAgqnCDC4eKZ+mFYjh9C6BGcIvvYVlrBk9LfhA2WC3XmWDeB5wivccZ/cXQjg8exvr7yn+2Hh
qzJSB37qYBkhpN3HlNsqaCdh0c3MSQRchUte28i6F12mLvufwzxoNc63jskzfW92zNaj5q6cDeJN
nTZkUpwacTacXMV4UKC/kmNMvJayCgD+kURTgzaU7vNQHU4V574VNO73xYVs+nwxTsuI9S/U20cs
DJgK1F8KLqSz2DR4ic+HXspwldOdqfXBL3YmnJJX5wTMbwlasYs3etbUSi39uNJNRV9CYbr6PkSf
fN98AsNCtFgp6mM2ZR1HCnf69p+kVus6dkN8Z/nhkmgx5E3O33FpAFk6pyECDj3G1sI2noGWdeVT
L2qidSulXBLm/2o2kXX40bLc1s1Xd7M3Ax+ayyAbHIW7S+u/yMQOyLfq3ULkq+cTBKBSoZ0xhG3I
4i6hBalMW3dUKhHAots2SnyBOs++mo+E8UVcRclFO6kNjEFdkpqIihqIed84LdXWBxHTe/+Wkf7S
ROYdRAy0YpzF5IFbDI7c7L4LfnmUskptv/kccuprAhUNjKeWtcV8WKEAnchu7UYz+OHnYnoGNJQx
Zom0oYWZg+73fWAxJI6SK5aiiQO8E9Ea8daiP1VtRWFPTp+sIxFuuZdn7xVoAdfVpuRA4wBDbCpp
cJMwww+ozbLZLdRKf7nCV1rilKxR3TPIo2DJs0DbqIDo0Y2pCdYiVU15Oj3nOS+6Am947eBMiBUS
D/colH9XVKCXYk8X/do8E7ZeUJUfP59/nAELhGaYAmVl/e21nelBEYGukB0NC/C6AWUIA/WB94Jb
Hnay2TDrmf/PMmrALW2/fHfv5TmSMvpfoHeOBFXrVMBylXWnMsiwGzYQS+Xy+xzDPgOpYptnCfWy
Fpo+iY3MhAPyALYIgVNvEDGco4NPieO6B8pcW9XybybbZVhNB+2ag/Mr6b8SGByj4QeXtvyB925q
ap76cPDVHyKKX/zargN8NjVXBtc+DZumHRkPnqTm4vLx8o4ZtWistdSPu+swO+bQxAv6qcPJixqn
Sn0Fp5FVa5EZf5HYudy4I1U5J7OA+P7VauvYtU0iCHpzbpu/A+axNXrvStix+u55dNsJY7t6tQ7v
0cCvMYXaa4Vt0wmIODTQlA/2jDxx8wI22WZ1hm1ywDk6sdcF23vR18cKgz4w/qjJ+5k/XrvSDkbi
fcJpxYynsWJkxvrUma3vbnOHGSjo6t9hjnyhZd1vR7oEmIG/A26gOjw2jTkLahZvmBUhq27+lCiU
CyMquy3kmU3nN+Ie2B0ZaRHdXGlfh/k/J6+cjA0uVQiiVxC2RxjjkVDZd5Pa4x/SxFueCQVTXw55
tWKphePC6SqMdUvjvV3yQE1be5okXm6b3/oAhgQIbnHfSEQEr2aEfq9Qk9EnCLLTDca+sTEeA0y3
Ge+uClbWHtX/llRNml3Qx+jzzovGlmqkZkirAEP4OlCzfQpSoFLe/+TV/A4tzBfydbeEJjqCFeKU
gWX1KI7eNkEkpc96hx1u6pD254u+CbjTNhKVbUZXWmUlMHUAq+M6jYSv0OaB7Yn3Kik1wRbliba+
ffCPmbhYMUiQTIJvdDEJRLvFObSa9ItO8wLinoFbbFlWgXvc8GbW8hCPhdDVWTIg03nLyMWWydfr
2jbaYnt0GUKOIAHQl/zVWHsmrLQBcJxSsKgX4M+LNhhYG4Uo1i+J3FIGwnlNnkDuHn/puqMR/NaT
VYZs3uFqOiHaO/r66DztLvMxKS8O7knAFBRAHeKJfMEJ3DX4jOg/9hGlxpM94fTfDRHjw0I42NUs
FHigAJf8Whqy3+xO2nqq7fAVrhWU+tfz4iOs6PrUnRkWntd1ZG+iJaS92cw5ZuhXGmyYY2CQB1LW
oM6Gv/F+BJxcJoJEXcH4DXLZK8TPGuoMma59G6UFI6fvDnsXbEIrhQf2p9VpsFX2wb5WHBjU326U
Qy7MRryJ8WVrsSJt3rZyLwxVFSeVsOjp80G/bhJiB7oVVcjzquS/FKOlBbSRlMhxP0/rdPoGpjZl
4T8Jp3wNzhKG7uurzmaDPOYmSt3cudUZ7XeRvBllYPyeXlC/gbO+WTrRMU/yq2Ii37DMd7Lr4PZ2
Gww+8rSMhNGp++Eo98CDUm2RmKiCESonPb2Kw/EFFEt61/7XjD23MVt11IAdYnFXIhqUdBClvuW0
4B8qv47Vc/fXs0uxbiQocG5DCKR34vg7i7kSUPngbZV5GGdjWqhQrZV+fKet6ZyFHAUSWlvuimgN
uPdcFnPCcC1eXK28iwdcZFOH4pNJE5U8bsegHNSb2JK6gWo69OwgQj7yp6mfZcX7bdW6wVIXmKeR
NdYsZKZK8mprNDpJxvPyiBV5knigdy2L1tVsSjuggJUMO8+RTFQf8VCeNlHwZvwQXBPwMnvm8reT
1BVsVb73dH6Moc2v3vFpPwTcmAyC9YxHzXGKvtFHNSMnmJ594MnSd2xMl0JOugJjAjRw/72CS0Wh
SPDufDnwptng86UGtJQ+/1XOz7fUZaaCnxrYcI7y1n8kkZn8/OsMql/ViQ1dB+xslfjMsiVVNvb3
FX5tGgiYMsN/kJG1CYS0STihy0F/raXLsmqDLbGp0ocJ81xOvv9IcE41TWcNOdDHSlMkLXVjoa8D
cVtDKm7emDL6iNIv8VYiAj4cW0aQUP9HqPfikq8p+DmJEMDZqUeZljXd4TdZ9TnGY+mstauxmo0O
VSNFzjga1Crb5TWZrX2uU4biGCspgOd6ptHZDlYOONmG/8arkkXih098cV20Hu1HIS5nEKwDN4xm
D+vEv1+8u+de1a/yiuQcWkkalsNdzzS6Q1htnWCMXx9PFwxOB/ypMX8nf9HZ8CMUvgaqORjIPcx1
nF52mefVUMzC1kq8QmsHNjJaVnThtOP1fOpt3agc3Cc3/DaFLJ2a/Qd3oRlspvkWYW1RdeQDCkwg
IWfrf+WcDZuOeD8MVLePjOYf8l4k+SpnVkjph+vnsNiUbCPTQQvPaDWS7poTHmJiRkE+h7yP9ELi
n1h5P6VJ5PzEmklpy5XCIOia1eaWkHUJOTkmZnSQ2Hf+EJmU4wpkQgiLn1v2q+lZs8xuFxyqEAb7
osQFZ5YzC93L7n6j8Tx+YNWmf2ByaU3YdDZA4FE2C5RSwrkBtY8o/xSPIzAQ4diPCPu4gYv0Ee5d
v5pslLktRf1/yGR41Ov56dEhf2liv4IIIb9da4mdKJ/kzmIYapWMI4/EMNY6YQNTlsylkipuNLfE
l1/K+TndpD9/O98hiaCRm8B+7Tu3U8iRzxpUbA49dYtoRtGNkYNCZdHXtUgZjOrA02R5bEfoxYJZ
JQ4L5ukmU28MoPXHAUiXfk62UID589ZC5G5ME2TGIf8aqN1KR9yp6PT38ZsqSgE232UJ104leRh5
cGSsKm9kpKu0AeLRWOZSVmGrGnzUOl+FMoT+w9cgEZwgDRfRUJhbbDqSxV1TpWiZZYqX3im1IZs+
xmiSFSRrAYiTSZ1oGNO8Yj3J6mPk5YyhTBLXBc7ZpwAeeD4c1zD7olggVS+FXP3XHP+LS0c6wEe1
d5PjBl+DrqoiVAb3qIWyVCNK7c0p0wIY+xaEs4Om5uH2wx95iBhsVtH4IAF9iBe0s2rif08sOoiO
MtvNmfad7CQy8fof9qZOLiA6rCzq4CHEHCvKzVnU+nHvBB/jUNb/k9xZZRTXMZGomvFSorb6WsVq
ttTCcovVWz7uUTVxbf5AZIyWfSsfIOcnlQdjaM4AGSus/JpXrg7UhJXiXjTK5HUxmSe0R0Njnal1
7NkSlI9fkLr7kpTTHOpsQfrc+iRetnmCwwHnK/vuriN48CiLRE9VW8M4xq5iDOp30XtAkS1p8fDq
vBLLktobHZe2RoXh4xVryTg+kSfAgy59024NS1QhPFl4f1VW1WvDecwYmJhaUTwKS4X6/7s8bqr8
/IUG4q16Gaptqnbr+09Qzr+cVz3NU02X3/7yy6t/vPTsuDyl61nlcGlSbmjgHIK0kpULjClxW8lu
9rWn1MvtzA9PYC7f2fJ6eN4nV8JzVUJ2XUcJD6/ufsoAaZYwSy2NBgsL8gjD7unBKb6RUttL+YfN
dD9GT+ZmhWlnQrqDwNVWo9uYHRNXnePEeq85Y+LfNSH05Rwjq1PoyaraNu3RibsX51yOgSomadKC
Yh1aeRsfQhufLtf4TTryw2QaoCGNiRp9Ridre90wM+MRz7gRfMbruZfUo82hIli64FZJjGEHMurC
nCN3tJQxUydhjNaSbdFqnuJ2bPPabckzlx2q/6oyzJL4yWGvojQb+lt5xZmSfP6pwKEtc+t4LGUE
xYdHwDawacKgsCOQm8c7tK0fWNKoPteJhfuSRMiWDXqxo7zbGr4VClSlNsp0bOGCtrF1vPzlc6Jo
Fyrn98/wZ/9FseTJhj0OuPjztuF57lGzWc+ryzhFSHsvCDGtNvQQUz/a29fp8uFbnaqx5ig5ZmCT
l2dpP95KszbO+qD8AEMz0hfKZ3RuUFuOU8xsSxs4U0EXUdQ2APs9AlcjDCkJm2n1bKlcK9mq37lr
ZdyOabmIrY6LwYp9msE8bardntqtlX8TFNtQl3vcfYk3D8W9trIpoaUx+TRB+nGJOxEWxK4LEj3b
MKtVJ/ikO9w9WHFyp+z0ic+ewTUkd5oaS5UL7FQgniwzLirtFk9LyaIqGJTLvFOIaWmNewoKrCwZ
XEdICnJ7JvY8A0wWVzV9CCdpbQO3kI5fOfFg75NYN10TAoMXVy5cSyvxdiwILML9qmMumjsIhMgU
xBdnBjmY7/j/r+kstS/tY/hZQN0iZLUeE48hZ8DcyHa3dLJ78wk1ngdOgei8QqjMKZeG/9UDDH+q
/UOUPmFS5oUWpVHmiMlKDedcDarh/nvz3+iwns0QMklpz2po6yekdnAVPRv7wzsFBDYTvoasgp6W
//JHWB4yiSAXJ35UVnOt+KmfJM/O5kYBt6nylcgbBJDVV834SMCAMFNoQW9hCSxzzhoWhMxKAKwx
5JOu+zGZxRFDls0h6B9fS3NmcqIp47exX8XxkDfbBnDbk2L5YL5pkIH3jmdVu2WCK4EkjjH6ZQHs
13a6RRHuU6cOW9/OJiGmm4geG434ZvkdICzdkFlQvF+lP/hSYoi/qeRsyAO9jUXxZ3fcQ3SuE1O3
wY8V3wzWVNFJZTkO4cR26Evc7QZmeIHu6UPmlGBavs3cNOxGaBemyVVBkYH+B9NEK9aIZeWKOaw+
l3PATOzwxNrRB7M0KWKAdYAVg/dC2WRhp27kAPwYc8I8U2E4qChIkwTmjISBg/ul1xyjXtyoYKWf
fMMrB9VPugpiZuJcK/j1ZEBq1UwXJEQu7fiMH4d6C/ud+YBwth8JTOfiDUWkDQLtneMGrv1aouaP
OqoCxwl89hFTIqlnVtYYCgM0OuLQrJWlEhjpwyTdNOG316tDSFl+R0CQFjTcb+ck9HOzhwTbQOg4
+1czagy4BLQoznBly9RyzlfsOfuotwWCzQuzeXoig9SIa8Bhk9i/C8F6an7Ho2E4nQlGQmjm34Fp
XudiZiBQ6ik+EltTbHGpLxThLmunMyVFbI0E9xVBbWqqQJnDbuaGFlnhPUenLLlQqt8lxcCWPbs1
VmV1tg63p9dG6j/pSAfnC0vZ150sc1SeP80K7M9pbDPqXEc+PtLGgQEnYn+TU36uamQlmG0hS0sh
dhEh1TQ6hk9nP7Ho0zfcKhcHsTTzCBNDVNPZPy2guUr55E6csVVI59OKU2HLSabpLmx+k4//fezu
zJYKgACuLSe4FPKmJNR5gCh4/l7DMfoSbraUAVDepx2WMYs2tABFUeKZmm2iLvPwHd+34/dYkNlX
5GIZw6vZ74scJZYajfRN+HQVilQWVcROClxOjT8ImpfwVrokO0BtS4QByTnYWzF8Ul12pFYO8OyN
8GTBIAxoqyLtsvDn7Vpqr0PM1lPRtLMXq2qYv8stYy0ODzEgIEp8OAU4p4PwZpVCg2Fi+KQBI34G
MYE6qeL4Seio+vXshzvtp4TEFHsVw4j9Q5ZCkp0GdutypAyfkPa2EMP96GoSucKY7av5bHphlhEO
BJItZoa0L+HG2h5MPhj/xOVDmlFdakksmZEZtpCEE05VBqmS1cpThvY3b7k78eKo17wnDtSFrq6i
x5lEWU56SzEs09fGq9qLqYSOXajkaNnZ4eOylHSGq6fVauUW1SEdDvpY1FGkRoDp4P/Jmv+g1/TH
GzDUTjG78NJoH5DzJO3a5AbWRorc++JCUCqrSPDCCk0vsThRSDlD8jUiByDKRuT8M7dYWQdKZBEo
dqOzfSReHWmT1iidM8o97sqKNIVRO/1UkZ+38sjLCCbW8ATRPiP9bqGNT1vVIr42YqaJUCpplfMG
KaSpWA4fdLhL2tzjGT6i6OrsY6s8/0W78FJbOyIXE6dg5Qivns10gfKrhPCZn33qd/aZZyhbwggf
hF9ghKgPfkUesEagJwqQETeoXxBIfcX6AgtWiaNnqZ0hzHRw9jdwkAOyeEWxRbP3ZFzY6JolyDjE
BLTXDDGpokEaB/C3x2XnebXpauXkvBO0PrFwJwej97R06v4+UmHCwj5Rn0lOpPUN1juXoZqd74+N
hq+LhYH9XBvsZckgNqe+ohaNxxiIUrcJug0ItL/ixVJR3tRpp0GfgeCFBW978pKvh5/AG096AGZh
lwh5kMwrIav3pGqyepzReDh3N+U3N9V6K6Lpk/BUfvFTrxrK6dxws+dgrAx7yAeQl/Sy/N0iIc8S
0YXHdElIvV6P9+J1WiA/bpOLZaeeyW2MHX9R/wabERJ2HPkP0eEbkaMhZW2pqoFEg/vCqWYMKpfw
gnU9mlx2T1maPFALUZMLvHmry6My2pcA1gS/VGNEYywM/hmTBtNvJNe3SxgBxCo5FwsXo1zVCZn+
nXQKUmmt9w1IsOwRT82kA3CVJWzQBIhetGh76yqWv1o1l0ZK6gOc+oymK6ESmgL0ktaKxXWIduAN
IUK8NAgzdLSR8xOy7sULPi12fbkqtzKoeDuWAHZPsNKw7p+m1PXxt0gPCAJP+RyMoiZEd/qRoa+I
SzYv6x5zoFL0G4VOTZLrfU0CcrALkRIXWnMyNK8z9kzMd/g7pQ1FnfhuhCJpOueMdJ1vi2sGUfOq
bo8rExg/sT2fQ8OUU2yguMTaPY68D3DxU6Pz9d3ue8QCy2tVMMjAtz6aUx7gs9z4ZYcWSYxlwRDQ
lxeDrXvXjVtVDXBQvhftrf/eHG7m9ECP73oJZIVsBONGbEmHYICSang2MXtFCtCft43xQn/q36xV
vGenBeAKZNWgogSEwGHIY59CF6j8vInp1d9byQSRk6eZ3s1SDKb8QE/fVNKjcb90hDZDoTa4lJ+O
R4ZK3RCvLkDH78Li/qQ/7d7zHrO5wnTUb73d35SlqR4LcrN3ETCez7cnfTM6tPuC3kEG9JkKuO/f
nwrPE2e6Iw67FyfdfBBvlVXnVMbvy1kKHe4aRqbqU1DBMfl8UH1+jaFBbR0xpBjfK9gWSicniQNG
+Se6rIQfoLn9IEMSrsORgadx/kHBy1MnwBHj3OaExOa9QcuWUCjEuSA5sI2ZkL6pKmPp4Ql12iZ8
E/10Epo9hINsLkTIBy3l6S16MLfcxm0+CjQrx2guyjssLfApObBMBslSlqcaO5zGdvU63WZVjD8p
EX66eRqHj3zZViEmUl0/qUY6d1iDUWZJwzrx52Yb6/6bDT/Fum0eaECtANPC8JMzrpWvVwyWBnvj
2a58h/LacB3pS/i2Ve/eV8bgA15V5jV6zWvoYpopVynW+vJTzmtaMj+YeUHFoFZdYJVrlJHUNTvU
pTMTzyjtDdo+gMkKCR8hAXRrooxwM+3DRTkijhn4iItFNEoPBe5gjqLK1swEV9Q03lQAn7hKQDd5
onb6a1KV8+lAgbLTxtp1tg+irpuURNU0NF5w8q7qvdc6di9ZdSIzruFzCdZqrcbdjJZmpFyIP+Qe
f9zj47/IfKXZO9xD+4rXtlI8hMeDqdttArtdbEWOAiML6wGFI9ZxWUNZHePX8AzVtemdu7UKM0Il
Q7LyUaS8fcHEtER5xvjm4edDpv8hBC+PsL4bNarnTeWxJlE0a8qXSUtaU1Xifbzyz8Gp196HpYOf
APiCPT0mqgvVwjdUREVN00dv11We/3Ls/s7JACr6CP0p3Qvo0O3NV5gsE8Ct/sGpQheYl1F8mbSJ
Hh6+bAsmKr58FNLGVYzVPmWnPkbEZrUV1xLPuoloa5XMUigsw3vQZ6wLdtbSeTQyABS19H4Ev2ee
FEFI5K5/c7xbe9FC2cCFJ6iDSQyCkqy0GS+0Fygtkw3scbx6j//FqLJQUw88uzkWdc2y3KNood1o
SJsTce1NGLxxTJXcg7P/mgq/W/xNvPWneZA5pQd0AFG+ChbhmlGBzB2pcj/2CRmcOPXGcDVDuyJs
aadRBcALLGjf6EZCRnZZKl+KutObfKNwwymLsf5yykh/+H0MgJaAkYmhXI7CmFYOdS7e8amSu8AA
1rsDZ88vYwht18gvOlvq/z4erhcmGwtZZwA2L9VHJK7W3Ouir2N5VU7TDNw7bFKa56lKtO4U4J52
REz8aTsIMnbt6V5Lw0eClDF4VeBi0s2UC95PXOCu2n3jSr1lePVVhLIK3lUz4cdzJfq+LfKkr/md
esfQ9+HXnrs8hgSGt1zchTvbkK/aBowdbV2Z603XSJ/+R7lHvMNjlVer6xoEfsUx6FEi7b2gRqro
b5hPPN1//eTSteCT4UzWPr7CceZqG0IjmoDOd1fSMCqlLcwGT4AWyVVUjIqV14iVTAcslJYt8wWV
kMrGXi1tl+Ke0v2VoU0Rayc4BZ/L85VHS8yCGCwqYm1e0Oic2XM7BJuewQWrgFf3qyuSchlSCKZm
OLO12PWi3EVEi5NLLaHuh2mwMeP3j8ssYuTL2utEMxQW6cmBCMjMW+UF/Vwqp4muKRTXFOjzGsza
ShUQTQ0iTZbe3s11aUdISK9KxTyU6b1OfmTax22/tfrhuCW+AfXwhss1qt3a7G8hVPruYvybuIfB
pLkr73nrMfIDyWzepBOMH9sgsZaKZQVzC0Gnj/8W/U5X/U4td7VU4oQ0jIib4DutdcSN9eime87g
ScfLiFvNKVWvTIfjuizqJSxQLf4NCgd5XxKb5NcPgym/JKgVucM3hyXRyVBaAPP7WjDNER88CAyv
68Pr0mMGQq0dobI0jVl7XYxL7XhD90MHYrZq6sQPoeYwPQLQuLoveqO9I9dHAIqbSlhvaUHRCxBi
0/26NF0OcNHRdXh1wUs5Pnge3er2su/IqJ5Wu2IBMZeEhok9NWbTbyyWM9QNsD+7Zzh5xJlHD3zL
GX/+Wv/fgcAwvQg8gomMPkKCnJMLBYE4X1yhIjjZrq1khGAFAXm/7V5T0DigYzi+TIw6jNGMfA02
/9yGju3e6SOLNjML2QfINpLKoKDkfIer0obPSGkeNUyXCmjUd6FpQUjwxsDXF9gxqvNQsAVZRO+J
r+xUPaP0rcIbaKAKYT3nef9qaSf6IyzsAxHOWmmQuvFQheJZqvoBD7RwfGPZholzYLxKS55nK5yC
eouSDw1f3a35HjP6gYsBAbROt1/8hZuoS3B3KOEgrP4JRIZ5FMyiF5fe1UYVjRhm8Md0+DjdmhkO
oTBevyr1yNQTXLkXBVhXBb33Yicr56jJQqp77pSzQSXmbljdXMtcTWw/kyBwz59HgFGpf02mw26R
+9kSS4OOshs4H2f+SFWw8vIz6cRnCPabQhwCHihCFMNeonnuEoZQ6AlaxIY3x3xEN4pKUczRWP2W
jZeQ3uZoo7Go6l2s2wJV9Ec6SGRmv4itR7xvmIJ/L8rrUs0NcFwuIH1AFdAuu4LPamIPpASLNhBl
ApzxNem2n59L4M6TEgWbYjG0zXuto4ZCG7h0hNBAyS4uX87gQ6HE06TgtyaJu3yeozsREqWbh/n3
dqEg5y+dqdOg7Cd+Y2/TUarbR697d7T7BmzQrSWsFW8j8ZDyzI/cEUEkfXmK2sZ6SLRfGvgWGrYr
n+CChdDHtdrIEjyHz8WlbWeWz1WJFq/g2/9HSUdtqNddDf4BjzRV+Ay7H0xrNiLIVFqQgnduhiit
4V8d2bgPXg1UO7/J0AH2SniFLMPvUFImUBYGdGL4LpbK93qslFQ23sIOz5x1Ip06EKUNInYEgrqL
PwP9r2ZYe5AZtiTKfFabSSI+ULnF9vWV/ywvUVYCSX1ADyksNn4bd5Tcm4yJC5F7j1p6mx7i4UrX
wB3eDlVLDLPfd+IxLokJTWEp9F5ywUgnE+0vDmApGj+gjstrmP8pEvYKDFC6b5cJ73azrq3ne90Z
Cyb9WcoEHFSPW/leViwNahhMjQsHMnvovpQPnW5zGbHOPIUi9xIboEg/XR9aXjJlpRWU16JlMzhn
/YQ4zSqAO2sQIt7SRE09gHcGrsevKU8xEBJd7a2Yz6smaYahp4SV/1xiLyQItUZ8k9TpDXxbir6f
rz72Fkt8K/oSHv2y89F7alB0aqXebj5Sn8uXPFNxhJCwJYHXZYBxm2CQ2DfvfGIj4HayZoobp2ha
e7LX0PWlg0jFGriHe9UvSkGHGisfgZ81B494WNMzNi/FH8rWH/9SB4taEUTVLIonZNvjtd3ueR9m
1rLrN5NWIIpz/5H0Zn1qPuxIVE/u6Izs68owBOIbfltmq8PYNOD1tXzP2NUJ8fAR1J0HuDnfuHAx
cK2XxAeHcqBQvyJbGEzuKPIJ2rEEl/qhjJAk0qwfC/ktPs1ZqNqAw/C4X5QBUGAkRsV/0hvjFjAY
yrUVp1IC6txDQnwmGdgbrCNzN3TmmNz7oizMVTCB9S7grHy6Mx9l6krIjcsZz9km28U6IYgrrsko
u+lheFpOttHv89hqspyMXeQ8A/v1GLyjQLrFYWC08UpEIm2MoMw7jCNOaQyCNw+vUEuFgWd2Xonl
21UeX9/610v7UcR+kEWLK1T0QgZ7GTmndLo2e5EXNgfvrVO4A/jmyfWHkPNPtm+cABYBnkXV6+lh
U0cDBvEZoaCpxavruFw9FujueqI2NP2RAAY9wz0TyN1JiIp+o9v23vTKeO2Z2ahb+nL287YJZlcC
gHAj5SZe6M8pAV6sps1HBw2+CIzKvQWp4QqYVe6Idoy0H1Eb7iYa7JPHylFfa3c2ILINmg1FYABt
5kkMhf2PMLEAROPyeDL4uI8X9rE8gTi+fa2h34J2Ei40ygCw9PuMBTgQFgxdKHFoQ2kOmdd+k/Cf
oQBq+b3w49ap7io9pkih/pQssjz/5dA7DTQfrkzYVyocbujdc5zkQxQyUbqRWDUqrEQ2zLU3n9Wi
GRFcqSeFZBGS/T6z0xicbUViuC/XA2wf81sil/xHb1IRGHOaWi0qCWtkNVSwGpvPdVuIyR9tahva
o43fWAAA1bXYoyyXIHj+4Ka2Vp6JU4pGIsdLPUEyBd1GMs7e/rnan7ZD2UFHrvZjJUrtBgSEvFax
kWjk62fmTnPE+F3552oJNHKnhxTIipbZOn6ve3W/jpiJ5Yu3r7FlIsF2wRbZvYbLm81PKM4krp6Q
UsjWt7FIikQIOy377h4yVOfM0BUmpmMXxZNjvjHJSGv/gr60ow8C/0vnjWkDAGlDTtyPJh/fDdxZ
cvgHwxW0bYzzL+GdRwSQPIHfm5DJWQ6CbdON2q0Co7/KmnUadmA2SMbJ+AC3q//QRIuDB21/G4wy
t0Gh5rqJLl3IOYzj1y7jrMCspTMFrXHxP5RdgQYQLY4gmfnwxlUFH0vIaBdt/XYvA3vW7CA5JBIr
Ui09rTP2lH/tkCq7T9YhoCLzcNjVofSDwRN10F7er8J9IF9Cbzl+jP3x/fHUCfbV/kc9L6Fdjovu
PbJ+waNq+mvglD54OOYqAjK8HiRrevlOdrkiJm/Dz59K2jec2VW0wiRdTDwgTCrye8NBgk0MhVH7
CQTVuqNokmCVIF62S0BpS6AYg0+AX5q4iiUr2Cb8BRBkf+BptmQdiJSZZ8Y/wjStxFO1hGuJJBds
jo8TemBFKggaEfP6P1GZwbgOynNeArp/KPYetnrGrwGCVTheniwG3tAvR+scOUt5FPloSPreQ0O5
Ik2zxgEa4UxGZXCDUovlORf56G6LjbTpN8edNKteNS75vD1Qg09CxcmIm8wn84W8ofK4saNJwHNC
tym7Oa5N3bowYrLR3SUkpGmvA+UJIwDG4oYoODKvZnod7gS8uQlU14a0uq3o9C5hA52RrToNoPhb
lttpKH6BNRPe6wlrunhvlFGhmksSoLADLuayztj8ydTFN2agFDxJ8u7o2kcCdwJbm7pGzB9rRdi4
wM0dY+QJzbkL8y2K/VYkDZfYHRkGf5722Rq+YmXuYgXLO9pwN+ryJqmDscMubH4fD8IarAJSX06y
k9ZooK47BgarcYyIsxk/WfxDyo2tgOpv73nv2vvsZ+ePpZ9Nka8j0jU1TkXQBdq4WyuQ1zofMr+i
VnhK0kUn2d4/tfvrx504ooHdXG+4rAS1p67ymTCkj8Efcj6JllRo4xKSDIKnhdX+8sfVfmYV/WiN
UvcjuqjR4jcJJjqbtLUHaV0Kika+jDzFTjsaCGYCnFp2BhQcHDXB7PpsYcqyXSvpYt3r/1Zfxs57
NGddbv3rln8qsyWqlwpnumCIWk1u8SZrdR/82y/JLtjMCK4yThCt/3XK5hGhPQZSKLGBuUkraF4v
CHm7ppR9TEvm6ZyZ4CDnmwPbfULXcujLnnWARKhGOJm2Yw8dvTZJivRGoDMN8UtrTPdoBZuUsb1q
QeTcLXLI04QdykJuTByUsMs6okVqGv658ZuH4c7wS7mledIVT+x8p/Rkypf4T0Sy8KypPs1P4W0B
BcZBx68fXDZ03cC20FQ17nezhpKQGe9Me4NGWCGOsr6mHdTlalv/a2qcEA71iRF9ZXeVBpFhnQsj
Y25MvV7NJ1BAUtOftrS2l74l3ttsUeCtS+Eq49FQVgLZEeCkC+BntMJ/+ioPZUjJSvB6KLEnlTHE
xcWeeO2PMoTsYwtrzmGHWsN5kd/vvbpB3lebZw4Aq/LSzwLnlr6l/cAfpDpf2/g0vc/cJAofyeS4
c6oIKOVofjGfT/awaovl1DqIYSrjUCTkJ7ctnwVloAONC/skou2IwxGSJl1gif85f9rl+oz36LUM
q6jsUeAH+vTbl+1sbMRll6J7S5ei8ELLNQgBOcvuAdE5Zzw6AGS+agFtPOkWTK4bG1VqOSYJl5OE
lPX9rpT1diYrF4t+NcpgMZelu7u0JReksXMC50cFJxGQBVHL1VN6GzztWFWiG3uo1M1llvX6+gpz
ihCs5MUHt89e3n1oGuYVv9ImDdshZbxIRbLnxbim5gx55laZrWIhfd/BUXToE4B03NT4h0ZDvS+S
2rk5HROnFWtCajd2PCm9xjkRGbRPexxZuR0z9EnRt9UKoc3uYNi8yCFlL3LE1pQxaz6qH4kpiMiM
LyR6467VsVCaSuuggIWK0+VfdUND6ZMkVtclVpPmVM56pXnqQi5ahAWgHLqJc9BfXEA5QpkL5LdK
jLiXD0N7WX4FyOvNcjBYf+WHWlcyD2cxdsOoJd9h8zP8GS4kLahfN18j4p0MTqVVfUTvxJSoRIpU
OFG3rMoLTBSTuZFRqELNElt/nrR2ieVwpcQjEpPYmVsMY4xffRiHnSVzj3NNYIEllLawudpMtO0T
yhEcu9p6iCW9zSnf1X32cq1kkipWRY4+fEboOjLHibc2cElBXTCvWQF4jY54/+84zJHIVBz6tj9s
eoI0QkiKapq5RFE7rfK2TMz6sb5Xzfdr6HSH9Dq4aYRsbRIWM92lZUo+FmHOCTw1vnK0BVFfpxua
RRvnG4A3t/k/rMdr6ApkaGFa4zrDfB1/1GOsgZX6dNaHTySEkoo8/IqA0i1cQMwex3o9rpshF8Om
UJw47fT+wkltkIka9fXLNJNqYEORAr9ypS1pkO/EuL7ZyMq10i9r4EMB0DXnJuwpZr3Ashfk5Hme
1A1qZEmERUbknNpJpRlPcdMCAormFKFZvPdpIHvoyJdc6fZGn5BYgxIpufo+lVhdbMgJqsGtYFGZ
bKSUFsV07EX51V+fxNWfRFSKhEXYModQHC0PA5Q6Cqf5ROns4pLhTeUwZ0P8GfQH5k3m2srOFGEB
OXQ/tmyrb6NagrIThjGHHwrlmKrUcQDB9+soCtws4IYIe3e4xBvKaZL7SWesWC1aTHTkepJTBPic
MEml5Hjisv2L5/1p65kN5uS0t7sF9HUuuEJOi9Z84FUbvTvZxkyEy7Ri4Sg9577ciZ0/O2yoZqPY
t/BquRMF07HsYrCaKIi2e0ARnKVKQPItjC0I5ts8WB/ArUkfW2VOKM67qVy263TrHeQDm/rop2Gq
C/1d7EAuqLe8DA5t/r6cFI9HGTA9yPvqjgw/F2aEwLO+4XM/F0i5ovwsa2gcF5P18EX5mFEOTeYo
4rpWdqbQxdWTUS6jBlzkv+RgxCU+UtzBTUKAZBSCg5Sy0IEcsNbTdIKTiMMYwsNarN8hVZEKal6W
VlcKFto2fyS1IzkyTt6uGanzAsUWk0Oi0DB1d8GG/CHXT3dzic3z6NaX5gfDl2NVNJwl9RwoYKzh
qfN64BX1EdkBGMur/u80a2tB6Aa9rhJT3i9BeYABQncypmgQeQ7O0k0ORZ6FWf0P2te4+xle0C64
xPM7J3Rdj5udeHqBrF9+tmc8re6FVh6ytfa/eo4sytE5ORk0x4ihhhaHdrc8gZ90qNOy2s3AQRUD
JEcs2KwbPAuIZu18J9/wIO12lv3Xng75tbNXKkjwWk1HcnmJk967gEqbrmkvJbdWX2V2PdcgNota
m0RzI5A5xdHCBhoQ3sbwjdOqDgrkIQvDtwUssFD6dqxyPImISCsCYyYMiyP/lNTKh0TzvIXxkxSr
7mpiMUYTCFzcMFdUX9zuHA10nJTKFOVkk21oGaTnQBOofvcNEmZGoKYzDCKVI73Mmbq1ZyAT/NO5
wjRsVMDGik6dkF8by2RQyvTKYl8gBbVRVDdcN99Q1EbrqoN1rqMUWJwaXvdvKNcjXFJzZPwts1rl
t7ZcdDs+EhGl+uyQXCuLuU9kfYMwT/sij5CfbweVDZFb5CzJZN6nqxDwErtpjQyFP5/c6LByFOGD
v8CEI/pYiusnQzWijWAWIv3WgSyRuJJ27RbwUHR0iwzWcdrKOqOkGvNhbRUZcUEhB6zJbD2y8ZDX
N+4t+Z4Q3FAT5IOZtUeK0kwo9pTwPiZmKocowiCdJhMU2rnB0p7hnuyomlOCFU26yYpcUIpSxF0R
+jR3RUUWEqtrVSIZIs7BE0WboJGE1HkgvnMH02mpPssjlwxP8By29/2wqujR3SSvOXd+5ZYCPqNj
Vnod4C6uqrFL1KMJSpJIZu7HN4dpE3JY1bVAWRENxy3NcM1T4/2w4JVqQsJnlxcwrRU2vIKV6bbp
cKNQvAb4Jj/YMNJm9OH+iSeW8bJOPWJ/Bz/yx2B1EMOa0Khn1qYzSM4c8FQKL1P9AQhiuldIIUHs
wumBrhuiwE9NOuMVCHfBlazbHlAbaxyBC6xKdGl+Ha6H2H4uXfMFTFj3W/y6s0xfW7aPG3CRNvKl
DWKnZvSy3vX1yRg/oXdMuj1tRzVVjo6yUI7mYBqil8lMiCzQZE66BYtgahP5Faf0kJ/1NnMprnaC
w0xjxX62y+lJ0a4nCK9nvF96lyksme4zcz7sPezsDfnvo1fanpEiaaHpBk2SWnLwXsM8+QkR5DC2
VxmzefTVuHxzw/54gOphjowXW+PY479PWVROHI0dDQCCW67rHelNoElPEP1bDvG+2T0aIaq9aluE
WXQavBngTd7tZ9GPwA82096Gu5z3Z9o0OqTQTSgUD0nmnDkDtzH1Hd4KpR+BIPOElc4+Z++EiK10
3kZMKOSGMN4f709Yri5kKqbITKNUe7JlSx0wE56RUNEuN1uHL5nggQBjx2u5qPVNno3drFcPjQ0G
ZgdKR8idy/O06x9kjftwdY7rmmzKpY//gKgcw0SBQuZdtHia3UUK/8YTeyEC2owFNdvZMSmGqNBB
+ejQjUwPRDaufloGKHzp1l1q2486Xfhgmaxl3kEUTTptqFGX5x3FCKVY5ZxHVvf7EikOGyR7WN01
/6oWjGwVZOvhlEDCCU8EUgKVdOKERuCXJuqycYpxOd6HoQchJYT3SMLULbaMbqpLsal5gILufd2T
SjSOcF8vPDOaqZ8FOWee2R+8PHmnt161QBklEf+PeXxvA1HIXxpP3dtexoK3QV9lN3uU0nlnLP6s
/8VsZdQG0o9ZBIJXr0ruLhLCXty/t+i99OqtvIHGyPaJvzU6SHB2hQDyt8Y64lXIqSCrKech61mD
zCpUwzhnHP6WpMSCaOZUqMlCaP2hvYILFhanUcNaGBHuLmbhwmezCQizar0qwdaEZue9J9KI5eFL
4nmDC361a4WsYGdjOjW3whttXykmEUZ/ESBY9WirZBFGXSfT7UfTXhQDXt9zqRi70EwNCL6UX0yZ
o9mP/eAVN0akrZROMvqaU01y68CtxRIeRh2Lcjt6KFoAp1XJgptqarUykozetpnjoznW4EoEJj+Y
98ahLT14+XNS2GHYoLeG2bc2+hGO1ikRobiOUL/WmDe3eId4gTHuRr/qfxF7GuesE4a5u+NHY7ec
kzMfwGI52WSY7P/EIoiD9kcCMwsQrBwdKOWAPyo8jRB8arJ1zjPJ+c9mxghgmirIqs1q3zHv/Nvx
Pl7PH+EWP1NxdePhK37kIVhgIupg2c2F998xF7t7dmASsYvoXc9W1Ec9dY3NMcWqUUwt6klBICt1
eY9LxVtF/dJBtteueD17DjF3AVPXEB7qL9ohhgPnoKn2WqLkIR6/cAvcGGsqFMdYPWyNk+yptJsU
47xSUER7PLJqDInjboFrg7X5QBF2pNl96TW4HFzkM6uaB34vVFm1iU8q+Y205gXD/vJEGPnkRBPY
OSPyuLsWJPQBD4esUqORYAXDG6NS5E4oe7YvU9MqTYQbDST5YqZUgBhjQDGj7+rSBRI097VelktC
d7AbOmTeSQrDBHLo+HF5Qeos8eldfKgZnUfem6oxNR3NCfQ1GDqUrndgfm7XOlgO3/XRG0+5z3Mq
B0Ahh8eZR0rO/oabSbfTDHt85ldVyh49UxHDvLacfx/MUkf4DDXvq0bN5PEZEm0A8Fa7ngQw5aUt
6Em1IEY8RXUn7TnwE6mCTNdD4ixvvdcFAZADJ9/Sfh0ZPtB3rAb8K2QMdA2tGRcRrnvzOXSxvueb
Yd2943DfbFJGhXv2mDlhesmSFQcyhQXFVh4oP3Qukb6lz2WOaqoAhEEjYshIluc51BKXhLMxDdIU
Bx/LW13tnn5uj8xKFmwSF3+ig80ZMIkveQnNIxe/SmkEblp3wGoPEa5QjOvdqtJI5Zj1VVCV7YRc
fHbOx2RZHmSmvpaRx5evv83/QXCagk0N+4M+Me7llBRBkiljGdoIFIt1UmHPBtauagp2rX6v0Ld+
TtA47U1XbmyuXNfOGBRH8fhMmTrAhlCBF1R2Q7HsbnTVbQmN0DZ6RrZiSkYt9wMdyMmbKiWJg4+o
PcIDpTlDoa0ws9m0kynCkukHr5rfzsycE2k6lJcUPMKWC9Iax9eoFfoWj8YLWfvL9eNmWS7I/E7y
EnHuxz5L7Vgd82LIUBUFNhYn9cdE8cCMllRxOGEjJHhNfdxLmgTBCUPdn+rMQPIaq/iS5l5pYlmz
NTFDj7qX9+Mhbz14dxo3yCw/FyXRE7Mp+DzhnPylWUAcZ/A2KWlV+fFjix9TgZaFPOSH8wkuBceP
Nq/W0SLsjXH/+k7ohkFOohLBTsTUaTop2JcmDXNCRjHb6/nVUB1HemGDhFXfEI33ujqd94pGOK9m
T2oBpxguV83WrH3vrF+Z8DoLcuFGPbEoJbIfBym5k/FrZjPdJXkVQLkybJhkJgxwCtv9E3Z5a5Bi
L8DQgcJMQ05Yr4hrC/ggH5q2lHX4ar8KncRcNN2XeGky0JkAhj7Gl0MKOZ4hwKsCw6XfHV7cSuZ3
uULnEUVy7ngpJQ+XnIyDvzJXMbt7iixzvDKfg54KbNm5QfK8m/W3mSFhoi2dUCmYptmnZL5auVv7
T9GMPCCF6teClbXdwHnC4f/qhFyRuOKVGnPHOpSr7ZPXdcwFg2YsuuBn4e0Q/QmVTELw4YrZvKBr
uSu8e3bigS5BRyBKhIIPv7f/EOArjhnqBHFoZC1F2w29YeNFY+PSF+kNh9C66sxFwWfBsFNXANWN
Hj0SxBH687USPH5sRkUuKjSaNDov4GVEtqDdEAGOneAWZH3nDsZAlRARgqMvbztTaIbrf8fRTMY3
DW2QYnb0QeE2I6OSbnK3cyFS6rrSKSe6o7OStyZQdOeyNOVs69xsQM61HrbdTNGywe64Rh0r1KIV
neLWN6I0zoccShGjRblMzoYfpLoXHU7d6W+MqjgnqkzJlBwmRA9W5EkfFCYLqYpDws3lF2YREhnk
WVzFgldMZiZ6WHxbkxdHmCv/QILyPftQy5gikTUBwEqXOwsJqh3MhPCefutYZ7jcYUpWFBt7eNQh
ZYMIaJwRCy93CsDAp0F8RDm1H0t0e6jrffm5jgza1g5z1L6vvJfmM9RX+elHInRWKvsb6lrs97qq
64Qvo3eSTV7agrsR+E67qK1nJ/+UHR6sq6PqswadI1sXtOgHgtceqMZkolvAO9IwhG1Cj2hUD+DH
vPhfWDliU5AtzrJ80Il1xenmbZDlBf4a4VQy60crPRT1Or1OYQ3XYjWjYQl0h1Z7SduHRCjJEBth
f3HiDrFtm5EHLJJDQRrZD2t9rgP2fSI6ozWXLlN7QHg9Y4GGXsGFTLSYR44+yu+MT1aiK6yMsfrs
C4nbKvSoZIOoYR3EQ1XNEDAcDAOUTuqLTDLbURVfG+W5k6QWzQGbXgLHLIcRhrEh0W1KsVmGGTou
gYJ2anoqeUz3TeZw0MY5q0G6SmWFaYz7pQBnr9Zp8Zj1KifUAD+C1wF6Tz+/05P8V6j4gbdeQ/IJ
64ta88BcsRbpl3REm1xt2aTS7hfzyHhhEFbPjwbd/MD1N7j+q4gYT4H6wsBcjuMc0aCMDxSrcvqY
oYosbusL68JoBrOJJhtQ41jdBnB9yk/U47xOUpsXrCi8LuR4J/FhcFIiN/GB1eckKstCSZPxVYAN
igdIDtGQV6f5FqaFmWEE3hx2JZYfTA9AMhJpqQsvKxvCGluFPCsDujxh4WP7uI/pfDHUD08aNAhC
/4HuYD7vO/szM3wdY9HCBZUQoblpXl0T1whlykfBtoLtrRUDe8lzmKGZT8HbHXtAcPcT917TydFO
2GCwgHpyWv2/VDH/R89BIeLrtpwGfLQ9d/1U87ddk9alW1vt+FrqGIAFneCSJ76qAw/g0Lt9bWzW
lJwwW7rUDQJoWc+T24nBsolNrLAs1S36F9Jc5O7M4zXut2dUf3Pv7/wUMRrPEZANXumtGmOMRP86
2y2V62kf9n7Z42lkNYv7gwxBVg2NcKb7CU4SJdPQftsMp8UIjBOKJEa1eC8YrJEmIGKVpzRUuyL0
E50huaFz1t2Ib/tNP2Rq6dHAJlpzuRe1Hq2yTplRTuRoZwBriasCDaDFYUZMIc4/VihKP2ZT9jGf
hKvjujAtmU5h7KsZ/5o5qgBBJN1jARZKjOYmfWbsa81u2aMaCLoMnGwKj6AP+5IseJBFZrpBsalP
eLL4zcUERD7gYi3Lf8X+Hd+2QVdILlVkS+qCQGWjib8ACV5u5lSXUfc9pLYIXt6dCOhrozxXCQyf
uXPzP8C3O8EU/iIVAUnWafqN0vWp+BdfqgnOqge6aZE9gHhbzivxDza9nJ9VniHO/Xb2cTgtTPbZ
kIL2A7m+LLVUQDQLmougbjz84i+lF5UFEe39lb9v6nyS4CH5K4ddCpvnhjzISCa5GjeKPm/dug3/
LFXD9SS64FXSBBaxIRIZ9hgNKu83YpwSULpTQStgx8c+2FHxX60G9aIuKAMeVIXkoRSqDdVCm2Qk
JiGXyA+BVI3S6Zn70NpaBHu51nMFllfAMZ3UoUqtfLL1tcw9EFhPej3obgx1IXJAp4o7u2RMl7vk
Mkdn1STdKSYujpVwq/BspOn5hNDCarX4/uQurkV+v/2OSFiQKzDLOK/LskDbiE3hs1r3Vr1AMjA0
7/KR02nyAXUE1N4D2a8zsVN+2PPUhsoL8UgV7ccQhxQWp0MWXkvimepPlNdlEOY+PaXuYDOVqlBy
Qw4rL8KebYLjKMi/Hl9t6EczN749tJaY+f3eJpsqyB7a8JhLRB+i7SB2KBiRQFDtBmBOZRfbBJLj
dtkto4hWR7TBkWLT30GARtjaDVDDcaqyg2+TzKxbgJDPQFXzjT3qjqxrW5rfKPCF6eSsksJb3azV
wJPHYROivEQBaWbfMfeLjndzlMGG2a/B3oRRUyrQBtxkc9fP+Kz1HCzL306cBVJDYZEdhQhzjHa9
uuUaIKFL8Mk2e8gd0CDHL8jJLUma2TFlUvbX8Q6My+YCAl5pEd1mjXbH7TBD6ZX48oeclFIIQcJx
6o78NSxmxyd0hpPsMB2bLZpKU+u4TbimvQS9N+qWOIqjLqciiU7bThKz7kkzroYRTbnli1B6Qg8q
NB1OI8dejwc4uo46tOTfWpBCjS6ccWaFUP/gugHKQ5VDrPz4EquX9LqF0kpvTubtlAJDPD1G6MI9
T0nvuu0cFKZBZrdSc5Z6cTaNGEmwunHRk5vYcIT2NPssSGTWZMiZ1YfternxYv3axRS+6hCJUfaS
Ihvfx+M2iU14Wz4M2fK7j7wQgYSjltN1bKhXT/vcUqHkTMOsrJhuwN9bUqOkG233BzBqfsp0TcdC
1APBGteokEgYOcwXfPRk10L1y1DDTOgSzg9JB8LP/k5R8Zz7EKidtanG+WgE/coMt42V/lgMaMhN
hVKO//Yd0MX0U3IzbM3VbVt36+n50AQU1/ZdRDgIfNK6kJcqHtg7Gty3LKHNTwuLn2l8mdmtWD+p
nbzEXEMt7jUDTDDa0TXKZGXKJFxBZQimIsQwWPW8Bvi7uCe/1xyg7Skwg/Qe42b6hSFSslFz0n7e
+DtKhYmdVpvDuxwVrr+HwXXa3BXDQyPFM8DXJ+NHGzyreswuZq3I2UUd5DkbN/acUgJRAUmcxUPa
bIA3ttl6/sxcqjjDHw4CiKprbby5ICoo9M8TmXTUpBzQZp2E/omaoq1MJgsuxRiZEciUsmAIsAH/
Go9UqATlNSsRG/wXYAEQf4VD8mLxohFVxMzPveWUMP9akAEdwGsCCwgv16Pn7NQvqVuNVy55y1kC
WRKwtTocixiXViT4GH8APiOVCmokCe5aqsznRyeB+nlM6wxB8i142bQhiJKMlelr5L0QBvS+TRcf
QcvX2wrFLuGoE2eQwPU234YSz8CBqPUKYsFGPifijyQE7+f57NE/HjgtsYftpj63T7p0IBeDGHSv
S2b26WhWW+Ofb5XFKHd+bRMkbOsn9Oeazo28keXdmFY+qkZAHAFRwpFzxuHkBXD+hqLowo90gII7
7tdoO43LMhZp3XFg5k5u2z7M01UjhKrFonRy7mPz507l7qVUSLoT5QVnryJkPjh6DQH47vvPCD2L
AhUsAa4q35QFa2yaeUpC1UeVa8IvKXN6ZR1niTLX9Za4Dv1uU1UogQFJXJSJZ5YF/tLMBixNSboD
0CE/7FFU+MuNME/E5J37+Oh4Ugf9S46Qv8fGCrqIQk75AkDTn2s9tzyaxun0OvMeCAmHJDXKIpAF
dDV4rqwpADmZdCMZh7BXjyxBSi17EkFYvdwKN+n42WoydS7hzuRsKaxJHHUqyF3VfFIVyfyDtx5Y
4LGae44ZG1rbyUGsPvZHvUYRnYdzdMZilNs0+khjpha48sKz3kdPgyyxji6YR1fwqoC3lA2oNQiW
C/NYSmeEV3lWASdKBwruxcqK6owl9a9ME131q3wid7GZuG8aboyr/byQdkRoigfcqybPb0ko6KLa
LupMTdusIWGJaCnwZdyQ5/+Mn+oajeCNqUESSopMfB9JX16V4BUhdLgPMWZHtHg201xDbfqq9Whv
uZcb4Ur1MsSLQnq5NFOix8mbjMmEvbX93CErBTFzqRb38Xh7FwQgurs0Ahh1ybMshHUcbw0t4i4+
ClasPt7oH99Fz6R242uR/nIqbrPCPJrglcawnSs6YDcS7ScC0I/hcTkhxEe9yaArmlPLOBfOdfGn
7SbMYFYb+3QQX4EqwInh0l3MFJVatmQIhLOvV8KLe1BPbPx5RjJ387Wb7VeCh5UM9BAsLBJFNLPV
r8151QQMKVcoD74JLUBJuhGjme6krAkwyJODfu9mnqdSS0sBt473S2ceFE2XN2eWxXPctujt4SUG
GHa2/7KhK7qgU2JFQoH/NTcupqdhtze3jvgxdPgZXu/cxZFUxgcXhUEhw8JzthbehmpUWTpKib21
gVyqxoqqhIMN+GZ9uUNsxDuEHQv96nLCHRaONIniVLixlOGjKhoebrNzYJkEg+6jcTbWOYS5wPRx
seceLdHx53cvwpBz9SFn7FY1yNM3EPItW8+BMEwhtP0mAaV9qCWuMwQbKt0Je8OgMI2AAd9NJOb8
gK6XcCEz5s5BbDPukSD0oX/QI4h32gfE/UhN56pYbVTI1J2VGlJ9se6qUMKzBBSers4+MVWLBcCm
dSRTjTwNIUiqJimNCBSyxtt0MTaimMgedqPVEsqTcONoWrBvMWeDCzPnlEAevKbEASKAoCOAh02W
tYPDrxc9l9LdesmWXgZ6ncvJBfo73rTAE4/9uFfftr+kvJfzrFUvlBtmoPqAXi807ndv5TFp4LV9
TG1pEv8eCUJKq/UWA2SRRmGJBRayG0Yum+0leZwzUacnmN5zH//kOohcoIyJC3URnaC2N3NtP6e1
hTa/XGOxcOBPzte8AZoZc9YMtsh7kr8no2F90/FB2/FCOFO9VktX0sGeV7AB4hexz+JUnML7gIDI
2wobJFErntNDrj4BmpEFPVutzrS3TS9Fs1u0g1Ri5yZEf/AhwolS4hizSTr6jh9yU7pF+FbKizSH
fOMPHLAFivHMifWhw2Sy2YFj7i3nL9O+dRNPnctWH5CyQMmy1yE/aHu3p7vGM1rPsuCK2luiZVjF
kbSDypPLWaWrQT0CtTgrpcp6SED5wYnyCbv+ONxy/MlCIr0nE72oJJQgo8JDej24rXcFHJExEAp2
Zgd+INihbtFGlHn2IeGtKCbWYJ4kVLbm2K4ZQqVnJ2CzCeWgK8l+4f5N19xTUXSeHqYDhy7YfDYs
Wg2Ju0caIFcqn0Xto2CWJUXvfEZ7Y/Wb5j1khtshtrU+GREPBuqu0ucxyGLOL5stqPkKkkThAGyd
59aLSZNLAByqgHIzAyt0ATUuBKywN3OGM9FzF73IlwjmbamB/8KyABEBTG5yAdsTZ36nMOkNXxXv
o4isL9uM6Vg1K1dzQxQhsh8KKvBKQtR+IfGX9Vh9L/aAB8nDn/fKjfmCRSwCNBIoM4+rcUd7AIj/
BfIBLFjIcgTfUykQ/xVmkmSREFgi99mZOw1TIFAW4RLQLMbBwWrVQ/YEg8EO/aPZokvQa8bNBZbC
yoUaEVmJqPy2exIKxaw+0T4ltUXpNLehkGFP5G+peL5k+rCqC+4D4mg0L5LRQn1iDUZISgPrTztc
PQbyRIRgJdzEw7y+9AKwC0q28Y5rPGW6rKUf4Ihlmx6aqzexzljx3HO2Fb0587t7szr32EkjteHW
oq1ZUVrC7ZOoobKbTiGhyon08c5nx2xx9I6tNTlSSpIDehBcDMCHNovqivfQdUIC1j/aPriakTFX
yU0kxD09tQUJ5DkLvnmEzLViT7YMEBf5GD2rdV2z1nEgtc6T1vaZa4hNpOoKzbUAICsa+ocy1VQq
S5JUX/nAT9cejgUYpuYD46N7Dt2nhNoQ/Dhlo3hFGqlui1HdKOGtBW/N6syRBsgZQlPYeROmhi+Q
Y0B6lvFdMogfN4eizi7vR5h1m6DuqDVObk2gPV6IBKOjHNTs6ucXa8xmVh6vCjVE7eaOVOHkoD50
7x/R52ZXSN7Nlj50rENXt1ydDXKpzSc0V9AT4Xd5w8njuktQ79zaLdVmbUyqCUEa8MaLrJmSfCtv
CrOgXH2tnOLl/9Mi/s+hskXlYFHqsHARDzyxOfWWRnfNciC9TBSn5Sg7sZO08FaNXWWt63xorwuM
vM/jqnvBJxRi9lAvprBpBfmaTiSniU9o2hOL3gJtCua2mlYvb370fi3yQT1fir3duS68t18E5dXb
wR29iiYnnVtGmZK+OgQA2vS9YDVLd20UB6ajc9HUAvDARxR/mjpxiIm/EYBamHNzVIXWUBSObST3
dwAJ69E9A/KnB6sSvmcbqMccH2PXIAxaaPdbxRFABHGKjcxzRAu7sUvT2M2Xks9HlnRancED1Osi
ehUDgwTSOwwrC7QL+e5s/SbdZodlX5ZC1g861UpxSJqKt7+aIwe7nVsD61GNWFU1Pdotod4+RDBk
JIIBaOcnJP6w+0Ds/alsa8KuQmQv5h6QYpGkv+HyQM7WR09HWxdERp6YEw5mL5+/LCTZPVo1DsOy
7szfSBtpoRmJwJ6WP7lg1w6yHFmvFJeTVXFTo7JMtAnQQW97qu4Lk0hd3EiTr5o/L/aT9Mm9TDAt
ga8YfaAjNJUyFE2c43bb0kZBjchRfs8AbjNprj2OhM+yxlvsOLnHkxQqFg41V73DvhYAudKksP8V
y/WwefyzXYjKvy7HpabaV7d1nTT/3xODQ1M0UG8Fv8yTVnmB+bzdxhI6fyNZ5/gqiZY1zQEZIcXI
FrVfDew+isJm3MnRV6jUsAXSMZRhRRJiL4XxT+rML+bPTZ8H/RWDzBEGJpD5QG8/lsfXov+GZBqL
SCHXeaq+EbGg7BDl3SQSt4JVAIJhLx/zlZtH3dwNSxhaKrsj06mns8N2+4E7F1mLidPkt9m2T6Gl
eQaerVtVuxiMV+mEZsF9MHUVIwbmZ9xM2t3u1J1i0thRBbvwZn+cvX/IN2YtW1tVqEzO4gEUmU/M
3Ygf0vX7KCtAsLXTZym234xuyna14mUHidIZfZ6G5cKAfUoBkVeZLV5toP/1T8VNPCNEeQvu20Wr
87Ug59zlWco5yQedgwO4EkOT7wf9zruvlzPauUYA2xLEJ2WOsKqTMkFF1h7T79yo2gHJIzsDg6yM
Qxb0ohbmsu/Hv7zDLadQrQhbVT1aioD/DCbRCHS4/9KXuwx8LwgbBxZrc4kOwNHBkSHABEZUun7O
Sqn1wyXt3dUm/lFgnuONi7IKs4rJZJLiLBB5E4wTjUFsPKXxCt3RCNR8IBVWj9scrXmr4EAk0Yph
ldYcoD3MxhH237yJ/6Y+Ml2N5wJnuLGOgN0Qoeer4psA0bBD5pUgK7AsvxlLOv7DZDhQAzdUbxVW
vX/H9UGaKakgTVRRjWoW1UFiH3C1Un20KmEUsoV0Q25pehHwc625XFdJvVX6x6Vb2qCdpdhpraMd
f9Cr7Lfr6Al1dm9gZWetdxowgcVADwz5r6y0QYXuypWKcasHEZRBs1h2pEV+vU5VYTZJ5l3iScda
5O3KiZCtFJmK0dCdrDx8fNgNTgU121jWeG9+LlCjrQF0kxBOrIIs/JMYyFFWtlM02zDhiG7Z49rq
mlt7k+60GiM/6jscT0XJIPCuYG9A0C/8Kv+4zKnJWtI47GY3spgo9PAbpyWoyE6YztAbkQusVsHd
mx9/b+eh+1ou+Zfl5Hp4d4wx9izWEww4vz+KPG+xCnEvghNFv1OLWhmzOL7uW5VRt6gTjJuPfRI/
g/8LS00rA/66c4/pkNDDJk1lggEx4P6gWW8nwAXEYqb//lcXHCTONvXy6o737tfG9AHopq6y3g1e
YLidH/zNu5YbPX17GURA+rlZRJ5ObzELN3kWvnOQERqJC3/xd2p6dzwU3AxR6doVY24kZSfzakfo
AtUwCr+y7/75L4/vdavepNiwG/W1PxrDIl5FiyzxWkOMcNww3nlWxEcRs++sdxnE6OjjXl+yH5VT
9DILUUpN1cZD/ZZ5KiM6+sI6suZL7GFRujzDFJsaIJjvewwoKssXoT27ICafukYMsGv/dvDsuv4L
WweGFhRgzXZoJHqm/zxWrWMihUpXoi4ATFJ3M6OiF7WKqnhVSXNqPbqQFKDwG4OMRunU8IiSbXVk
YnzJ220qhKrNRX8A+1hUutnPLIMzSxkDhtgDilZ0wiLdoaZ6zmZ0fNsxV+lkrdOmNriV8/NroJxP
5RvmqQsQU/7Uy7D/XKfWNXvOfSkUHUREM++g2xKXvHJHSydj+ETtMKlIdXgVAnF3KU+NrJrZo6EJ
0iaWx4avg3NK6jk1h3DyjAwRXwyCDVPvStdFb5+0C28ZPei1MygwK19GLllkDvlXEkhr7Rq6l2SR
B0yLZ/kK2cjeKpsJ16LGlUXj/liAxHaPZyzqhbBaRZSVP/bCggU3EVUlCLrMf1iv+269D6jJv7LA
4uoN0pLEreDCbvU8qAQ9K2pb3UIJywW0Xox6zIe5ikyegeNTAdbjRqeDHZGvkHp+ZllHF8ySJsNP
9rP+28k4FuJEkGNrDBNAKKP/AJpkYLmStQH2N5lxfk2TGGARkm/plHoU1UK2rFlKNuJ44WI9PatB
rGlMByC/U3ckBxhxU/OaueDR7VNih19NU8LwJQMpZXl2bb7YESaYBJxR3SK6OhQYNLtiEaau57lu
Xr+x1jsWq6hYjjDGi+BJc9D3KIZPZC0Giyae4u6bmTYVUqjR+MUrFN4bGlVI5MiEwFFygq/OYjOw
DAPjxPTTTB/36WdXg8RQ5uLW5u1wNR/VwWVeSZZpyjc63mFp1Iu2Rxddhhih0VapAmldBB9qMZFR
UwWGSxaazcLFx42IfgiT+NG4H2QuLfMQEO4RmgtxtR42K0FLu2eRI4PTfTHkkZf3XVcZZha25lcQ
RLT7rlL+sxElfZ4ADnqc6WyRGP2h/8w8w2blfw9VpQDChxz8WOxIKjl12SxlQJU4CzTZDEeiXzEl
RBIS1qLwP/tBoQQvcvxeIcmdY28zq0MZ4K/kmRz7oDakU2xWGesG+em+xxrWAHhvi5EO9zvLjan/
zX5sdHpkAaPqVSE9NAPRxUMMBy8d0Gz8OnN3wBx/RIVGZWIO0nSKdyqlSfK7JsY/vaSAuatRwpKI
QlK4gRDXA/jdjgSOKJzfDovrxp/1vqyi9itVRnVUrNdKwaMvZtG5g40HAxm4OElS2+TdaH+yujJj
bAQhM5XEjnuC6fb2RvVUUelajzkEEPRyDlOSb/ymUBNziVWqthscv56qd9Hxo3wzPr+FheeKLSr4
Fg1xuA5zLGTnFU9bpUAIrW9kipISQLWLJtWUzf2ns9VeoNtm5+rBd61FnMw1gRnhkfULni8szwSg
Bg2CEDkcCZfwbik2DKDkvXrV5tDntX7R4Kuh8xRh9eReHfpNgXsdb6PBYiSBvOQsquM/SWdPUASm
u4myWk39jzjmhaUMYQe11WcDaBh1tSQu9tPsr+JZAiQWlebUhAn0SjiFcpprhsMiFe75y7ySkSmZ
KMP/s0ezYIcbl2EiEVCAwBJjr7RYj/QERN474a97IkpJQwgYBZdh5/parMyRBiG01jV30BY+46hA
WfXIrhF/xEa+7NRaQlV2oMobl3pn1WuwIJLCMqLHEYJqtnSt/LcTO75C+AVhvmcWfABkAURYnWP0
EsBn39OcFJFbJhjRN15cQba8GrWR2jYJOb6TxTFtDPYP1f3Y9gFG7nA/c3PNpj5cPuVrBXu7rrFy
hPASLHQZbvTlekCEbGakNA4nxrZmmQ/MEeDxw+GQbCW8Ky9o0jmMRYUAyF3a9LWEHHHapONi3woU
lwgw9voK5ZORsdYACRIR90jD5ho1zaZyEDkbEcNtdBLLYsZr/SA8wlStX27RzQPGNgVflyD6V68j
XmE5HpNOyfHlo9U8MpFtItRum3RAtdTNY4vb+vgl2h7+/B6/Ep1v5PhvaIKqUriQ9/s4Xb4L9vra
AjJORjD5lN8YqMyzNxzOVUxCw4Au7oWeDEAVl1TD5Y7Je6NqEkecn5LZBG2A2L80bWET9bVm9EVM
GKD8NiHONKzvlpTNBUK8zOKNEYjEg5oeh9iyywnfos+xAh+6mUT6KeCmstPYlpyCv8QGU8h5iszA
OWAMkWzFtqPRRYTPut/zsGfcBx4dHS/fYyTxQVsCVBT5mAUyV17snmxMTH/9FExfhAcGy+JJ4GNW
Kos+ujjKY6Hishay2+YX2Gchn6h6vE7HvfOwwwkI4ruVLv+qdMrnqpCnoIqfzKjBb1187beaFMg4
VVuVLykUEb80+JiW0qmn6TPRswmMTmvZD0tzvsT10bwsoSugWG34ZMpPFck69WbunnM/i/aTKnlK
oi8UFVNEXB3WM2dt0OYxk9RDC0VvclsjRC08RtViewjm7YhzB7xTLnv54wJSbc9YyaRu/BBtr8b0
hPMtq1rrJEHqZad8db2JZ4BlNmaedjEZukjdlIYX7bTzNrkM7A7ryA1P4GykQuvSDoQ2xyBx862R
2A/spyd063L8ckr8hjxVCt7gFRVzD71tM6v9PWAj+qZkKOfT1l42Dx3aqflcFSvdNOIR4xuzxa2e
C6jtFMIAE0fHY6G8olefKiOTSeKJ6mPY+zXY35R7kCrEw15VCVSO92yqOE3dSJt7SyvUqKvcgLNg
5HOLPnUeQCy3D71+AxsuO447NXj0WZsAoMOXvxr9+cPMmGUrXnscqwNvAW2GEqVkcA+nllkEAC5V
V2mRo/OroPtEugT0Z1TEpb96g67638JisjCgz0srOgGxRVGiwkMM5uF9Pg30WYCUhrvbrRlqmcNM
TkrIIH4x84cqeY06BrI/rCuRMAQSgO1hFrwh7u720MpCA2edhDhbul9PHYmCwU7td53ndTrohYXI
vFgaZp93NU8b1d73gpygfI7OMydxVgksf6ICjN2mXdLYuXgmi+KGz60dNmTY3eIn1RfzfxcoDjKy
r7AW3xVvK3SHUFOth8ZSocNipwWvEvvqyBJpG5RG2x8YF+/O2QqxQjkLEL79g9eSVs587w3p7hOy
OoOKi7NUoKo/XxVxlUoHdmp3fz1lct6dfd4qspAOx7j1uZ7GgwadK81pefrd1ulL/FwUEJif+Muy
9jPzD15n9Z9REyMJ6GEYpO5FfDqr9a1rwO+b2iH02wb51DVaeFjr44gSNCsSsRbmgX6dLtIySwpR
whIo3IfOqcHN/OKEERPpFUZigrKptJgkB1fGNADZRGW1JSR8UPGj0rkgNjAbeSX408Fzj9M+caX8
nXqHRRtn/CLoB6JN9be1XfoJi22pFVwfdz6RWLwqeE44fMQncbB7+5g1kKgrntEVvtqkdJmx1IF8
MNY+Qb0MM4KQeAOQuffmL660bjAP8Ms7gKIisywh0e3Rnjk3/bpTMmAmjmUzgBaQImxkL9cXMued
ImZj21vY837GhLhG+GVt7msKPOwpXEdhSDgOHCNGPbDQo+s3Qx/VQwqqhoOLMQpUwBeykinxkAeb
pPA4lqw3gFUKGvEIh0unNkcWWKtUI7BkSZcG4L/Xn8B0XGTZBhaBLtksrPoGLzifpVzj0ma9/Fdz
bbGPAOSQqYK46zcMJqQtNU8fQB/l9JzjDOp+Xcpeex3SM6MwUWniLh055qxxdB8yaHgE7vfHZRqa
I//pK3KkBCF1LjpgxGD7WrAj755WhyMRQIAHOimdfxQHBobDAXV277vQ2Fc5TmTDlHCSY7IqV/oQ
WlfUt5XzDaPJNN/tBGlEFIK8HGYdaiS9kvdiw0b2wvth2eKd3JnVf2MPj9FEvsyRpjvCnSW+vgiZ
lrDjfR9QPd9vDsoXBlvJgLCQI1PQ2a9obCECdfe/Pn03A14MwqKNkCQfcUbUHkFdTIxteMhKMoFi
kjK9CqNIwP2VwbfJEJ9a1d49ZLKzSs2b7AYflGbxzdmred2eoIlqWl0/oY6+BPttW67raAarCn/3
P+Jty/XQNcS9noqmDWozHSYaZYwlbEwUJobBEglipJDk+6zbD3JsMDhwwgo0oKxJP+xrDMBlNvt8
PTagvxPX0jA3JOkm0wCRtFWfF84IHONsbdHrK9n2kDqnF3M9W/AGMjc8kfCQ5elLpwBsubOWyDfx
FYhojwiFhRVSfr5U2goSZin985Uo7g9OL75Ti6esGaFtr0ImqqmdLmdDl9G98ewOte3/x0v3eM6S
dRT33BbnW99YsJqMTzXXs8vKowgXfDFe7MmJNIBw3ZKBdkXiSTy3MIKy6aBh1vq+tYgcyzOCaxtf
m5CnEBSCDDG2B4DIgFG9ud3rfy3wX7RpaXl83C5fF+pCYc5mJIhYLohrGvmBCYT+yR3PS/c58rHy
v2eOKZ06LjqT8uuwOIZNk0oW5jWUlsgt4cnRm9NbPLhNwJqldSstr1LPtXr5b/4y9mACLlaLe/PK
m3Vk5pKYpjWNpQc0Z0Za3OHLse60vNm4pvZRIh+f8BhJ7N1eMgJZMipjCAE65le1WkjLXUk14qbB
7Cx9dsGRIpLYWAFsyhJ9tlDbE8k1ZRj/pfZY0tvj8y3xRiUao+Tz8RMb7rUgsfffMuzyUv4K3tvK
IhKAWsqWtKNkwk7zqAiSOMmC+NBUyOh6sJt+GWJ9ypqaRtc4SRPUiUyfYCV+f9qHVprccEhglRoi
PlnhPwz5AGP0OY6CRk1/xeTJ7vwOS3UcfP9ok04+Mmn7JqdYXyZZ+0D3cHh3j58s7ih9sJ9dRFRb
Ygcy6NVuGkJyqLkDpQKGZJO4m/l24IJlNG0rBZqOV2uf40qagBToAgjhKlXYuyQ+ruwTw1BzxouA
CETLpM7jTnrby2KnIfTKAxd+JNeyaFlOG2cfNFxyaG2JMphT3a/AOvEpmO598quZ+SHOdZl9eaot
dS25x350OwPiKJD8HzO/mBXbnKQ2W8UWCwjfhrUUvJvlZHVuI57+6gGoZPBsjVJF1JTIBWrdaooS
Jps6Do1+UUQNxkJZN9ABIDsDKraqheYz/lVU6/GtQZffxXONJRI8qa3j35qX+30IlGmae3qa8PuT
ijogb0wyAmpnayRgWLSZSQhctH8fMOmdVlp9v0rbKavGQ9utcoPFx2U31CbPrzzY1F9dCV1v741m
8VnY9jlJdDlGkwhx8HN/4yaeXfY9fwoQneF5ZSNsYS62kMj7gx9zDl/eZ99PB2ImkkyC4RybLkio
+fWvpUxz60DLO07IbX2ruYlplbPWDAn4Nzqc4AP9b14YgWl4xWGBAvoKp+wBbr5zjTq+/7Zl6jLN
bsr8ULKpW0hXlkiuRiNWmoRLlwT0erbqXvF/28/4XN8sV+F1Eqmr2+IKdrOqseHrAI15lP1o1tBM
UL/o9LZJX/0Gq9VHjQIsW/jk4Sy6r2QXX+8AlrBQblT2ULlEwaTx48F/wAn9Se9JUqqRriqMORci
gPcReY5tU+tj8P4OfBDw1lZaKzVRbXMsGFt1JRBCFJ9MDOQYFDvxdOeVhIAgIxtGO6Lti337OVKj
R5MWkfK6WT4iPmQ1ogz34Z5zDoE3Z1tbP7jft5mhTINq77lHBioH+ltfc2o17PHtQihWDw8yMtE+
ctKayhXRfnyzk8hEg6TplrHF5gUco3D6utnSRTJ6In1sCx3cg93IVeM167C1fuiAfrWXh1oof3sk
AiSg+sFtUBH3hTAIG8qZO9rqAqE4REAAlbkIOlaCfw3yp/f+EB89BUDMClgAMsmT8khZKJso0WhU
3NTfEDSDwaWB6UQuBeTJEw49PAAn9oFdzDaKkA/BY8+7FfA0hLJatK9cXBbHNicYegdMnBhrVKa2
8q6yLWjNMX+h6HHo/Zhn1fSLSmLVlJFdgvfq7YjfDh4HKR0ldTs0DjFaV73sWsqM+8Re1C+sju50
jk+NT4leOBAgTSUOnDqQPbYxfH87FoEpt0L1a8r2XRLP6lcWgtIQ2iCDnWQoNqG0ZtKUYejoppDI
oWhZQoRCJJtGJiqK7S0Yu/aFVOxY/Ta/xzx/pnS/pYtR6tLBEa697MVXZMjmWvkS6+aii5ic/OPT
haFOWNcxe7LqhDax7E5DFJ/oYb9Hz4g3gTwHJxT29uMKH7WWNKC/vYVMGEf9s6hfkj4l7e2xmXFN
LOp59Cod3fYG5Cut0OAj46Jm4G+Nv0XK6sBfxodneKJxiryoJ0EHN+gL/j4d23HJwFkFVUBAl0gu
tsws+7cb7RXVWNew62YMH+M+EqHdZQySzIwjsR56YWUL2rU9hdZtRudY6v071eg956XPeLMKTmAz
d4/JeCWedOqQCKe45b0IOfYf8imPjVHFpYzeBwOwayWfB7xLAnfYMVpQqm7/r0x9f8FyG/jSMjjL
Gca1iJdEmwrAXD8ggtL05n2pL/ZcackALsf1q4/5/dxNmimgfDklQU3jHEL1AC1uKlvv3Evz7yNm
nsYXdItAQSmNeBZmdSgsbKFpvGdUiwUHTAHJXB5o0SsRQQLatN9o0g6PoSYm248DP2DE8gV0DiaA
jER0IOAPH10rG8kzqP1kQvBqHGmQxNk/OSbdYQ+lGtX6tJGGUhY2aIpuOfXDj7SuODhSCAMuOssS
nklEyvTpoWbyOqruS/Ca8a0zF+mWcZgWOeM9w1InoaRq6n8LzFwoR8g1HES01fWwC91X1tah/TYZ
PLR7cZr0XR07B+Um8hGB1bIW7EV4Ag705oikortOkwT1IH6KCKpLsREqkSwOrY81pZXslwhANlQT
kgRqrbycBtOSe/kyjWakstPqgVRUQGUJRewZVqn1QFb4rE3in3/j1Nb6JnMMip+HE19a3KJb0QL9
H/FjwVtETBf51ftFuq/BWCYGL165k+YoVsS3HG3krQ8pbM/j2lYXW6gILPVfLMP56Q8yXnXzbtly
/3kcWufzeAQaRZ8dSqyN2VxvtltPL9L/30WdNslOWRO2eRsGDwv6OK5hojxdnUyTdrKX3hAJlbFB
PLkoeQHFmF0ZYxkMcmyv+PLf4cezIDdU/4pyksw1stzzu+BPwgRHgqQBS0TBz159aoKeEuNN4Snp
mvKM43biSdKSGCLnoFRlMAJ/ddE9upO9cEG9sfaS+HDSUBGhFAXycaBcbQ8j0BH8USFw7YrpZ92K
T6pku/c4cMA8FA3egdI32ybo54yH1jzPbpQmixPn4Uouc69k+0eXz3iW5pzXDTXHV5JqWlIUq4ad
qAcqwYRu9NzfUIItEEaon111rLihC2XEGiM52WnJiv99k0OL0G3oPH14/CLLLerKHFKutMkZ4my7
PmbC2B6Q5pNJ8ifWrTph7X6/d5Mqkifq7AXRHNbPxl399HzmuGPkHsgtfxQnmnYoORUKQbqvGbVf
EnUD+mGP+k7+CdNOpb9jNrxL/KbyRuzaZwnlF/SKr+EkP6CbN7MQIG2IM0oBPU2rKl1uXS8gwfww
kIaCob12beJYUAqcXupYOyFC3H4T+1PVs/ghWCVIgJsBe/0GCZgQidjgI+TGjOz9pklzolENFVdg
NnsErNeCEFSe/baMM3bItMIzwOrlPL4Pwg/465KDF/kxZr89+Cig7dFpuwgtSpA8ce28bcKuo0VU
21ELP/cKCsfPHqHJ9pRF4V9mzoDME3grTDrNEpBTpJB5Fhy5irSLYh5MdVbVJIbj1hOsjZDEaHXs
KCT35viKPWq1TFX7PE1Yk3SCJTTh2VhLmqu2RRZe/x9CQDv/McfcIPKLHnkcbwCc33pXWqtXg3YY
QELjBR9Wr3ynYkJivSGl/mXzQUQaULPS0PoWELxQCxkIhyJEXbu4KJjyUm2fJDSce/KyLc8qQ9Lh
y//iqR4BFRXGOarcotEWx6olsVkEDj8Si07PpJ1yAqg13+arXV6j34uQCX7jRfEfEwNAk0kLt32Y
yrIvao2bpA9C8jYck4fCU3BXMCS+Gx2Q+7j6pcYynXXtNtLLOGstxJS+owxU4YG+s6JDtyfBVaf0
Lm47ZMS63Hz0kcyVLSdZSTb+XpbT4JDXk3ZpV2P5fMGbF5E8f4IHOc5zix6jS6KI3F8YzISuHvwJ
jAwJOPv40SZEoG7kdCOlsRSBa+NXTBNeLiodoaSv5GEpAUH77UnYJz1iRNXWwmDsck5RHKWNkHug
KoPCXT0hctD7hM1p1JPYfYCkC9bGIndkbTWCVLREP2COmxOP7Z7SdLPxDeaSYAHhOFjhexGskhwb
mujd+Y6C0Vgx/aqyaN800+fd7gVgu/QZIvxROYCwWj8C+r8w1aTaQpPVGG3/ZePI9ZQ8eK9JkX7E
uEtA+zR5XJ1RMbRSrMpMVjRcI2T19F23GSSlYHDkuAaXd3//M4iEn1nfVirOY20vfDzfcRdDAk0K
k4NHAWPbiWyOkAn+G0Bln6926j2U/XvL5wKpSndkSjKDcY8NVfrVwlNFBnRigHLqyx1Z413Hkv4I
orEvXKtWxP30CRxS0aEWwuZYxAWwGCvomSm7DhAkCwBJ3ISal+vlLeU6nLkMFRZqbDtYJcXVT7T1
VEpsVRJ3QsJztJKh4Fxs/pb6KRcrUibgeNByHhS7E8ME9tDAJkKBorTJcfiV+WIHOzYbJhGlbfp/
Qulbmw+hdA6pnh17HQyDLHhpvI6S2+/cocfTSH/XNoTgkGEdVACcrClsZghzvLUHYiLkB/kpD1dh
MA92DpwjdPU06M79fRPRs7aSQ0MrszIPfB6/6YqI5ffWwnXFneMN5pQO6Fj9yuSS44aQfWnLAlhr
sPb1etwqPiYjvlxeTaKYeQ2pJ6DAfSKmIqxfdodGkWwONXNL7YD3L1IREQnOCPIoJXGWaAerrrMO
GQP2tz1y2M6+df0T2CMTKAweQsONKOhaeRNOVTLK3nDYqg608+L+BuP5ip9kYVDIqnHioHpgW3Dy
cMfxnhYfPEE4/fecesls7jQcf2fGq18J2pX5yZEn1tYyxofyVtQEAy8Mz6BYeRDzl1nJjaGBzZKj
WN4HWCaR3Ybytf7SrQclRwUycJwhXV0+2d4fOujr3X7s6Y14nKxYYmhuDHg2tNNNBUJ4PQD5SccY
BwBzsb5g6/iCQJ8MrEYCSARoPhJimNWoratZWdjCVqEwQePARllF0dFgMH8lyjRwV5LE7MkY4uoG
veVYDyqKPezc7kG/Gqlz6Uz/usW2UeXaMW2+7NfBC6Ol5S3tAZsZSK36i4YPM+dTSrzvjgdInATK
rY1hz4naiNuWL5YnsY/w1HDFKNVdey15janxbTNisuxsSjGdNfP6pyT31aBJZ+mSV/KJVYuzeHbQ
Rl3t0/4NOPLjLx01C60UwzpmEN4LqHb+VsmxaqcntrRjuVYFdV4D3hBgw12IgDrgSsSGCMz4+Vgp
it0GODFexllp/sZhWLIxpFC3GX3HLvhnjVvgpiNdW1m+RuP3sKgeuiqQbC8JsriOYYgMAc6g9h3W
RXMvcD27FZPrdDQIJYprj3AvbPmbORwCq8PctKfvqiVksK6SIg1lB3uuh2dGTtqu8vbcsEAy+1Pr
3cu5QUMJoF9IvQ8aRFa0MnfcsNOKGIb6P4d67VFSeE9LLAd5VSBMJu2ennSjFVDHSS8Ryq4SmUXZ
V6TWOCvSd8ZWC1UK4VaHYxtNwEqDnBMN02C35HPw/nlbSXyGFuS16fQam0iJ6GZfcRsTNWzUyeRA
ZpTQc15BXgl2HGdE3XZliKYOWh5/7jRn965QgMWUUTEBrIMsIbOsf9jJEIfvneAPgQNvhxl/zQRG
mV6PhL8JY7LZk5gyhyrSf3ckwcHyzXNCThg53bZE48Yp0O8LAyau8vq31imHnJFsG4i0h2rSS0eL
kOcDMPFVwPwzFYLhCIOfvgN20OlYhGm9F2lWGBjcBrnJEG/CqJKxVzbWIvXSYeA/l2lTGqp6EXEb
rAqhjPt7SAupp8YMwEkrgXLCcDH3f/tHOaeE5QH4J15LkB019iRABi3f/Jtj4lFGbwPD3udEPxfM
H6mOxuVOBFmviheZjIHUIh8XUrzf8HVvkxjuYwfQCZjfuhzDJffZo9ER+edr/7nUegVdUuo8lQ5t
t2ot8VLKebn+lUyaO3Nd2LmyJIW1mbIm+wg/rLrnYUgUEvunEgZSaNi36ocQ0mdMmqk77uvF04/X
71KbEzU9ZaPlM7rY+UPmW680PyEzc+Sqm9kLj/btMMZkQyIMk3WksjmxMMyIxO5q4S9KKNFa7d+S
7h16q/p1kxHqoInV14SoUQJfMRwA+fa69gYO8ljliAoDEIlQYjgx2zEJEzQ6M87W2YFH9b2oNFsp
JAbBD2j9/HgA6tC23YwJZdTmwJKQjsFO1N2VlMiwvlg8B+ZqHefhqcjiKqc5vektQb8PtIVRv1/x
799mxRvsI45ChpZa4gpx42O/nYonahqXoMald3abpObcMwCYUkoIpNmx+d5c7mcRamTQmpRJEapK
ZwH1oMV8NC3ObI755U8rQCcSPRRm+Z/BVRXf2+YbkNGiCm3Iv1MbG8fv1dJoSgPeQbcyneUL8tXt
q8+vCK9wW6kQJHf+gjYWIl82ZpIrVgKP0OJiKUDIJfuUVFFiUqw+wBZr+UXBCDi6c1jiHkdv8NV/
tKm0t+q8K7FDMKo5n+OMHOWZ/j/t2oiZL08UHiOMQnoBo9hCa6dQmjbY3b6AupnSi1J7PUF/Cch2
EGyquMPyt8qI/VHXsAWVmMwJO2QdyqeyegWfX988I709OAP5MXwaWSfdExpZU0ujofFmebqAmsf1
YAdh3R8NO1744yzKFzdozS+zvCszmIYL6lmwEzuLxmpdvjWl9+wAncScvpDSamGihel4ixC20qG8
tdRtjOoO2f0hJR8WlL6lasAhUxMCOUiwzW0/Njam5loDCC3LA04Nsi73DNCDZYAGZmj33/krU4MP
CrEcBhW9iP8G6LDbTpd4A2BPmh1PLXY/S8P2P0JrsJ+1e6weu89HmjTdyxIZ6Yx2nfi0bkhCeV+O
5KzjRnJ5Ku8GfnV17t/lxEMUlZABBMj3rrk+ydvQSt3Y4xCEMkd7PCDS1JTRLySqPXYcPTzcm4Kr
IwkNbDKGKlxqFfqr24lKj6nwXawTsG5efltLrgFAt/nCQnWa1MgnlmagfdgoyoYhUfViQtdfhfyO
Civ5ibZ9l1rGlmyPEyhAbiE/1ySqDeUCpKRPFRMylnoheFp9g+HDsPODyFodb1x/g5CgJHSXgdmE
O+LQ2U+VJlxwjnVGtgmkrnVYWLRSkFfkB3tvIMHYdk3uPFknQC/UmMwcPj1317L/VIQX0IxdzkMk
gNXNvOdPHorv4JUq3AHqwhro0LPurAmVHcqGdBVl5wXuKaKL1UbvXKVlBK8jfAUuvqfZgvoGGV51
fSq55z6eACMUZJ5J5tIBCxywMb3GZWFzHrliOD68Iw0mHxjlPZrwfytw66ngy0rs24Cu0UdQxX0m
f1GmYIhjBiNTOld6f5WoqCZ4z/yEJiF5iOJlboi/OmLsyRLD29dypQna3VbjCKlWpkTyh3p0bkeU
zj+b8SyJkaQ4r2UMX/wP4hSkPq3ZdqsOhGFNxxQT+1HwbaNkJV3axEs3LF3B/5dORQjUOTcOIvUm
2VBXqVv38YHdia3lEK0Hz72wzDmS28WJOllF2QTMgulCDLF66CVWlb/x/ezJwZrqObylvT7P9+oh
o3qOMxDUpqHd7raBtw0cnr0gMsKsEbNroqNLkfkQhARkbv1l8eQlPoumKUsQp2Z4jj/gjPNMjQ51
n919xiGPfTpP0DdzZjJW+ShGluslLE/dUijme7ApfpkDr2m51oXlJoW0EIc7WgHNzHnuEzInKLbx
ijKX3feFahgB/9Uy7oyPpu/ThBrr9NSFBJmz4aRVnys61queiy+ccU4/+dy0/Py4nT+qSOX/po27
eWfF37udqKpuo/TZ6cYpcg3Yz89nHS8yXnLeq2RLrze5Qe8GYdGziKcRM6x2ANGgbdAe68iA5nbN
wbRYO7pHCf7z6npIdh+Qoya4dKz0GVTW0C+OVzK5IaYwmHv8ro8joVYA4q9vaOywcJLqvlQ2VylS
HZ+UpOtctkSvDWigzZTGMc+D3xsIESKzEhyg/LZAhMXHbaiYD6tOpZ5Q3perJBCzmr5pMyQoqN3r
kCdHe3unraWuUHZluojgS3RkcL+OlQ53AGIg1BW/442IAwNMJbxxLXt1wM8eUUkoU6f7p+Ae95kb
+Pl4R6c9Mci5Qzsk4ml860BbXJYNlajnvhP60+KmZJwh47KZIjSPPoWqjhdMgAR2I0YgZf5Rv3Fp
rThAhSAvunc0UZyqXtw1fGqV7Vu+5PZE3QK3mdZBXB90uxHkj+0K4ntybDRe/rJK0imoYknoR5XT
4+3tMeMKYQa/95xveiHp0uoBciYGMb62IT0FpYY85RoTeG5Fig4pV55HiEISP540FpOABvXZ8e5h
WXMIF8Ap9ZMNzELMKXYjcEe1qa4IwIg7iyKFRGn8Rgxuo0igSnjvSRtDGRrCNWIh1F4boyngH8z0
2o8H/r99orHlp0goz4ZJPY1QkfS1D4w8fPdyL2zagD2MFg08n0PwaRemwsQtHA14KIpwwAakUfr1
kVBUH+Sl5tuMaTWsc7YZkJqkXgoWbX003qR/yVt4q0B57ocRIvntFCmgXMzTYW2TYwlvO8xR2Eym
VYewv+ZmdXua1LW/W30IPr5YLiHE1rszy0ZJNEld3ONiYwxNlCKgSfiSPSWvo9d2t/AkQ6xgqALF
K9XS8HxDWFrxhCFb/LDW2wKK3gT0i4Cm51kaVc1+rzEg/36dhpL5eHfGRYq5eaxaea7b7obcZ5k3
/UnTBSi0giqQKemacNTX4gp7XzAlLAnSeZL+JFLT+GagO/JxzFhyn3E60n1snTL8yh4HrmupLN4h
iNi6bJ0SvE/8dSl9u/QjPB3F6HyLOQnTlp3dAphJnTpJvJNvEFamw+SswmffIdPLmE52k2TYULIi
A58o8YWghS4K2SfypKz2x6MGlnRltGRcjKN952cu6nOUuUjMi6hbc1hA0sBgwwrBYC59xvchs4sh
7W539oK2dT0H1vgDQwkIap5jr/KFVuzfeFfyTCVKTA7zu+1mDkw3PQN54giQMAXlC6I8E4E3D72+
qZNjvD9pz1eH/30QwjeTId+z3G/oxsFkP2D1yXrGTdNEDCrJOkFCRh1HBKbwTNFrvzMltsnuQ4u5
k8TyJMtneOOHrIMYLWfVZ2tmDxUXWnpIPmLyFIJoDCbe+hP1zE6UcOa39g4isvydP8xZHaXq11aA
YK3GdN4ZIovSVzdnIwrcxNm0H1EKwzIM52YkT5cFmf4A24Nmr7Zl+1z2ACftPD0lEjrjkw7+eOH8
nHyNcED8HTTSx5M3XOZxLbdbNISgL2yFGqAvun0YH7989IsWUec8SwtXtI2r8oV1bMUabYnIQjv3
S67CDGwIe6hOz2khJudVTi/QGbAQG3nVE25TlYvG+lTGQKWdLIlm5BlZZzJy5dTQPkZ61y2+R66F
3hxnzZI3ysTOEh1lPXuIHbUx67McOdAl0lXndxSuXele2KtbTUT55wU8Bpaq4crzQh/lMKYeV8+U
NWR2YdBAVgfsKY3x1+mvzBmJ/OSj6+GFGolQdQGkkEnImZgJwGR/B3EZrf2rTiY+6o0m9Wd/JHmF
l1n+wzqjfyV94x3KEHtZjAU2EsW+0w3jaD8cfALvrnIp9dWctHSnklNMMuOLf6ch62DukTKXx9Hd
1Iz49TTl2FbKCG4P6jeNaxvvAu85k6ETI9dj6S4yNfjDgvk4hNKtZ0LxJbuQqoBlFffB4ldvZgpF
0IQ+AMpEu6uApYGac66GSQLLkQlz/Qy7WPjVpz5aZ6UF3XXe9R6J9fC3/n63+bJg9aTeTcPDfC8X
fENtwnyX8EVccdiGg193CfuhgA3SKcWuefAR2N3pb2k673Cqg+rYsA0rhw1rVuUtK7BzjIYXnlXJ
A5IQyOyZmdXQ7ytOJKDnJtDDWjashxdP4lnr0pExa4sqYW2fMRf/MziknKN1fEU3qBMeQYhF9Dv7
d5qSfUa29u6kMqS56F4LcjSclRtgQOU2pKuksOW0yfQQmvxwv9wI+9iK063tjmoXQCLUvaUJImaw
AZdAjaISwcUsaihUEk/zVLJNu0mlaGAnk+edHHAwXbjvMpSY7vTV0WVLmoMEsQydzbHiSbF2TQUz
8432BKXLY6+RmCf+b8bMRrgMuAouDXqCW8/45gRoGH+NOX9F0ksg+TFWXYmb6Ucu8p9WPL8YbgC4
lG1UpnyKuXK7RcCtuTMGEVsYjeLKYNzismHHZ2uMUTnZ6oJNzTIg91cTsBVYZlb4ZjtkxAknSRO2
9U0XmJGnE6FXSvoPxuig6exloU5xi1m3MIxHAr/L/ccli8QfmPgCu8MF4Pk2etY5VOmJjW7xAPVS
zQn+GQbqPhMQ/lFmauRE0V6HG5q8pPtcGlR3KeMV+gP6eBYMO6JRexY0dhphZF8nSqtMGJGeb8DF
U87I0HqLs8Uq0ZEvlw6Mjqia24JIDGsiqFhkxvhPQcSwzOOpSEo15X65zXUihg/ng79pPnv6f+fr
Zjn/OsFykIrNZ7KEzDinR5YPojEqqiamcSHhpLvpLLHnj6qWK8uP2fVNoUyqwixlWTBMj9l6KDYZ
nOI1lZVE1GjVQEdRR0igL9ZDQfFEVqPYdXk9Tjk/K7pcIoo29Lf9nyvw6tmZqLLu3j6TxDgHmhoa
ctUH5nj/IKCRMQNblufFOmIya9onYqp3i+X3kPCY9+BvN97dqQVTW4L98kOzYbW4EZqatE0Etnxn
+vI3mHJT/reWu3cuI8TIbj9XKua+UQAlgOC03TFBDSGCshoYl+s21iAmLYqcBbZdHUSQfmiKS9jt
9LzrEJZxnFy02ZLpCtfHYjhzPMwM9WsgginyoHHPtXq1oquSGAJWoCFRtPCv23H6Pm6qwv3GoNHo
SyUs/xbf3mKQaHoBlO39+3RUugDJetMyCwWKyG2RyVkic7jbY6rVoUgwDKm0ojgXnT0XdkBYCIa2
RjVh05hV0aBJ7xT3JBqaB6UodH/Te1NwIFWakV53HqwONYz2/xk+Jz6j9vkQC9Z/l8TfEqQpRV4Z
tB0NKllIxk6tx0uHWi7wZV/d47gBYW3FPwrSZkgZAHavB6r9h1Cw8+VqmC+alNkwspFKZQUv6bFp
5OkY8WkjL3Eezl9B42vNpD0/9/K2eLH078PV2IfRScwjSvf8E5MR5waNf3SvGu0ulXlWlko06rVm
zb2L2fEVDbAzcr7e3mCaL1bmlfKJXVxfaMjI2EL33a//lcoLQzlKWYMPvdyIVsVmgWC6elzJtqeU
r/NheNy5kyTSthVJxXsr78kf9csFs1rkcU8JnPxNKdNCgm+WU0H/G7Z2n7sI6XwS78xmpa4DBadH
1kCm7amOkid/BSXZynNoqrhP+k+NEtu9QrcOfxwi0UvqbQKzmibv3f8/UaJDYNo2dktiG2v1sfjy
N6KRc50h0Caj6tvXZps7tTruf/NoHU8FsOHCJ/SqDHs2lyXN/1789s++bE9QpNOW7G/a3xtL5XKG
UpUhb/X8QV3FZEFZUq6QHYj+KwrX3+OB/IsvkBdXaYV9VFi8yT54FKFN0m1VkM/IWYD5HXlLGQga
oJaYvwvJEsxkgmMis/j3Y5xGYF5jRRdFLK3O9LnevlvcXaVdBFe8Z2QMzAJjkJ1IXCYAfiRHbUKt
Ag+Z+jecVj1fQ8Sv9IERU+CzcNcbmPLmS9tcyfpqI2pT/9fY8UlLgowJAGu14HnJwGOhH1Hpw2Dp
lo2RNDvNYGhMlRuB7kvyWRrVgGy6xioclnKShKyLNSw7nMpn0pLEEKXG56uB9hu7u1RXwpKDTB3E
FFZAjxXwymGsnFRkpBoSSEx2Hu9wTlycSdzhANHYk2q16fnJ4RLRL395STx1cRXaCkDsZO0O1gHf
CpZ5hgcqayDsOVDiG8e6FeVOwpxJrchkYnGEbciw/gQtM6zYubI0CQN1tdHtOEIa8nG/gREBBleO
vJ6jAHuSpW+CEz20kJBSmzUYckIJBvne3F2SEtb+EgDvZ9HQpztUFUlPyH/xL8QjDQ69FKAqsGhf
9aIr08jGNeaFQC92W9LYqLcKCzhKnPjVD342PTrgWjBhWJq3/LPOIDLhHPGcyPAs1LJRDulTukX6
7kC5nvetxxkZ6Q5yIViemavPYitCynVaYlm6QtSluXfse33N5HebwAeC7hthqqHAw+HEAU0Ygx1e
seivvGwSyICDeT1GGqGxDbe2O/bAMNRe38AQhgam65c6EsI4Rh5zA4/lWTe9NQPZbAfgZ1XJce90
DiN3L0c48u3JYkPoB1Nneg/ZIYCYXaN0XTIcoRqaYHCGVOcZh516cApbUUOWwVR9hko9nx58E5S/
2iBjtmZQ8C+gUOVO2nd4rSmflhL++L0cabDjTaUXtMDDwtex3wTueAOPxHmX96NFITO3RyCXpjS/
VeHlUwQCLLgvt9xOG6yWujy3ZjSega6J8mR1WPgh8DLTRjGCJxlYz9aHm1uCHmxaf15OR8nSdpJI
vrhY1kEdJb7Rkt8f/YIadARsBAMUqquRgr5Rxi1xpfx4Wayt1xLoRA5S/GM8oIuw8TJVTwcOyfZH
NQnP1t+YRGP/RZSneTzvMnYXva8EInw8HPmenzGJ5fkTkDYVk4+Q/p9b1ZHMcojcSaQb8kKTQxsd
RLoAdNC+XLKyNgdhHUMDZIObs+k5OY0QIH8dv4dxijTLm3ibNJSeA2T6i3Lr8K6PBX1kaIcyWg6o
eSNf/n1Rgb/+ak8rLVcdVYWe4OfUbsZfUtTdGeCJSZ+2NatOrPPJKnZtlx7Bs0SsJEfjGugy0fIp
unvhxtYmkCacL1/KOHKmQNIdpfAmVX4myJC/pFvYxBwU+I2GxmEj465arKGO3MYlRq+ZliJ4ILwA
OIEQw3NCwQHhIpigPekAsx8oyDXX4/uVnpLKuMgwxT6UehHd2/RqCwhK6fQgDLfI3uOiu9HDt/yt
/hnp8teVODuL2BeaK3Vwg8XePyC9qrQUFc6TfVZBKkMSBDhA6MAuNoGcKv4Sk6IxbgA4iS3TwD9K
B+JVB3dCLER586xTI6f/dG8cLc+SsXwU/nyJkf9fovk7PIoA0chjZfPAz+BMsfZNPyJDJSI6GxOe
jEwUdwpVqE5dGomAIecI9ROClYe4zS7JMZ+kwocXVPvCqeEloX7qQDj14Qi8GjqhZFVgJPmUEiwo
bgndULCG7sd3cdXROl+eFErmNdE3LyFt9fcJkeuzGTLHcR+OhtORB+T8wyAyMcvDPU8n+D6JRnlY
S2HyeRnMPLecMUHxREkxQtB8ovPwepLbsUr+COGshJQjJ7FlZu7V44m7kfo2Zu3CMiTpA2p/DU28
fkl96Yq5Cygwp5DGwCYxG0orDlnruu8ZAVu4N71GvVWX9ikzsGnDZKY7ioVXmcgHKQ1YDXXM22pK
FBdakOL3NWzk7Ce/8+P2wesdZ4BBvLFpXI/bHZjXM/Gu0x4zvXpRfk/f0qFDcum7n7jrIa5NyFtp
itoCuZ084PORO5raVwcXIqeh4CXPOGCVMdakM8pFD0DVE/Ahr+wO7FRbh/Qpbdg3oUaCHXaTNQsP
nLB6Md1tPmvS+BUPK5wXRyGB32CwJg0gR4HLtVkYYtyfR4vHAyzP4koJVur0m4ThI0hDYgrioRNg
HasiR0d2NLLZbul1Cbs2m1AxS93lSauq8n3Ub9tJ0reiZAhXBzjoGvhNZy4bfr/1KwfFdVxa7/AU
bzY6DBieYWfhdoh1bauR0ORCqFk3rw8YFKr5hB/vgv5qF0fDin1jFEkG0xffAtLbNkRCm2g8b2UJ
F0WH1OClOzZJvsyd1wbVay1bFE6mvStC7SbVKDUeoZtufXtvRnzGn0uBWkpYRgTvxEAiKfIjWZ13
unCCebVvCyYnyrGZMV/N29vKLZGJP86fg5q5M/aM2VcsukeiNF+jSfMQCOoATwf8w8zop9102yYA
18/VnUN+IcnBLdsinjb/zK8XDcu2tvijhbLXNuodGmpEswKzrIU1f+Nnfi6MqMi1yTi6cjrbx8q2
nCXNy9ndXZtkhzFyl/aM6CPffSjKCnEMx3bVsoPGCPtiq4zbiu5WopjmVDJe2u2DpFQCSgNoX3Zq
4+v0lSSllGi92AhWE8iWvxSZHF3Zbo/ECI8nZBhMSUPtKrLLntxIQcvlfcQ/3mBY6fVnbYifv6yV
+0BU6ucrtODueQkKlKT6s8i8AYVKE0kjdkC952ixr2Mc4xOkZUQzyxf7w1OcovVY9SSoyz2GiSrQ
4cVephzcMr0FxVDY9RmnuBxn3gHLF45VsJ0LnWAKLRB/CG2oOmkJFQCfc2NXOA/T0u37M53YfRkP
/C4ZXBrffVh9WuSe/nm4auj9Pwet1I5OPJVlp5ukxD/EZVjfgF3gBBpeHh6vythCxnNXoKyRlx4Q
AAHT1Sn3i5oLRhERcBepoCrKdPY4OSJRmbY0wsX5y/GMK5/FjA5W+jvTeiovN/lY9dzwQRt+WNRB
niflSYcVhejjnBTFXwQX1G5q6FncIwPzbOTaZR4cbuyXZYnY4E3fLN+CwleYeqRuZXtLMSFi7vIK
ARjMc528WDyjMC77e25ot66U7fBSnyqpDN2AqVc5MThOEgrOAOcG7TaYk2s+TL0mdDHTpusX5cDi
+dnTaKbRaQcJghz1f9SigekI7GUEV+Greog3UFoiUN2wWw6Fnub+Oclzdjb1ZLVIo6t+KK9zanQt
wlUCEJj1btYKfkE178r8pUuSMJfNWMc0OJcgU3H4sxQijyGFZabRN9VsY/IKjFJxKpYPIMfGQz79
+WOrrxZQnQOOoN2rfWMqyh54RRWUGALnoDcKUihZqNb73KkBilEsVONWpM/SREiCtFUoXgouukAg
24hDiF+5fUigVbasfsJvCZZGqIkb9EhbY+U6LKfZVzqn3OL74ofBQz5oNSXv23N5xv8mHW5+U8zk
e9A/iFcXy1wvk1m1BYtHnyhRwy/o06I0TufDGHRXDab+vVqDd4Fk5x+tt7V55/7M2KyOWShHhCIO
L8Ruw6xqdgnx4L9mwvFiW8X4EUVwbFWh2qShp0mgKGg8Jct+C90UD17/Dmo6qx68jh0tcJw+oMl/
GHirbFHAcO3LQxDFHOEMNtqV/gnk19H9nDcRysrrw9Wd+NKkVyVYZA3KP+BUd8hwPPqMbkixxjfy
NCMve8pWT5Zx3iuI179RyBAQE+0yfS8+oPliqUumvUIlbpdliPpxGZ6Fnqcy+xE7QsqYXtvLRgLO
kifcRqjkUWH0Di/Wjc+hWb5G1Ib+ytejRrNvk76WEm1bD8vTz/kaTlEFCnwJ6hRn99b3qE4x2kJ9
SSAhvp6uMsMLR6dnmSklCJDgTzOpHpkxZwz59/BT0yUkjRwnbnbmmBJKyy3hCZC5nf/CiWA5PzgG
4ckQz7bzqT7zsMy4GEqIaaf3znmp3C2aDw5rKZciGH/2KdO/xPpSFUJ6I3uZLGSo8vCwJi5Vrzjs
p0FW20vZplbcuNZKno7hUUevCkVSN1li0f2LNKM3TXAYKmOOFvGYUgLkJ3ZN873q1AtyJ0yLpmOc
JejKPaamNRX7ZGkPZ8Ub4CIVVMufWoD6QV5jxNpHXKizbayfwU4Zd6h9viM6sssrJG+md7DzgpX8
ReMOHc53YmXa5dSfWQ8dZDshJr796x0y1Q3HMyCWrnMW+u/CDHa7A5F+zIIUGZ8Lvy52AUr5lfWE
9LEO8llf7ynAE/pHggyEAJgwquoMSyqXzLeUmzVjCkL1pl+DjIHAL1w11Jkb4e94gieCAFmQcVTf
1h2rcnKbBwKK7KVX3xfwQw6omjucf83uC3WCtrq3CtoLSjtsb5Vr6MO+cpEcat7MXn/mKGaD/t9S
0fBrrLI/sLh4NdDBzPMr1M195ZG9h6t3UF5SKlOaYjroxat9A56A2u0+9A76TytPJgJMLY5tKJdd
ytdFAdnfIGqKp9+m+gizuGLC4pGOrreb4ztM9ZThdqPgdhb8lNQdmvKlT8SDLMFJaPJxJyEZ1b8U
u/m1v9tR2/Qx4BZ9ocaRKxJe6vObvdmuK6yq/Qr80rZKn3vzvlb53qTvzAr2QptCWFP6XC1BrXqd
1i46xnhtxzisd6AGHSJkmqy/zJjwjavqyH8rNgpLZh2gqORtRcpeW0IXo4bWpEoLNIh7Y6F+PJar
G6MLBSfuN6130RARQikSOleF8hKrLKSTakPPEpigxx/lTPmyzHiPB7CMcKePN1BukSkLQ3OPZfJz
C/e9s7zGbDJL2IRUsSWxkYU2MtCCL85bLbYn6HAECIrg+3PIz6/S4uBzFxuKa9qsOAXuZ7ZTH1sC
oPDFS5M4dxWSi1A9jhXWKTA8QbMBZE81H00TvrjBAWtO+/+bTUHX5yaDZ4QKHVGqNraXy22Fm9Fq
HoLYgKN+H18WnRZwtV26DXwGx+NvOWVI3ES2hlHNIKQ5WFFkQBvK4nGP3qHp+TzVw9voqdo9lZFv
1R4OjsN5g2LaQPuha2/gBqy+1bvLhR09z62RbK1WYoRvTJuMxhX+jpicfFcnvJ/8ecWYHQgvRdqf
oPp/StWbHWt9enB7E8eQ7sF1YNz03Mknz0d45N7xS340a89GEFC0Cal3l58vcf76ebUMM88S755R
YC7DB1YC/cie4tNvQVgTkfV+83vp4pLxzFZCFrnAjT/g0K+wh1LQHjJRvY4Vfwzk9cWk90QWAIjK
80vvEq9oqHMuNQbIE7O+xlDuS7rlhGSDqtpgx447a1WwN1tpZuT8Pmeca8A/2vhpCzLQ88aSOafV
wd/3+0EDpv0yXZgLTSvYbR4W9iDzgUOzrr66MLgcjaDsi2AVZoeuQONzMy8nbGhb+SGXegQHGqPt
39wTg5jWSyhi6pvYijCgndMyO7a0iWrIPg+PnRj1PGzL0OxcY6u3gw1Kha/hQfZ2tbbSyDmle8TW
fgodxLX59eBeGlh9hdDwpCARI+XMn+VI3YF8D35ULD77fGUz8fkRzoACU1vEn3YtjZMbx7ssbaEk
B3Mmnev0fccxWPTlEdxCDqg5AQ4bkUE+sPP1kDSPGrO40z3SSC1z9PxnmXHpwaItEB477r6kyV7m
ubaBnRKPJs1WCH0V33mMnaras/E3W+k28YQ+jsjhtQIyLD3w9+9ogNszATY36s2y8TN+qkVD7jhW
uXGVhQDwoWwPPxz1Ebxv7l9FRkK4gM5MnbkZJBCjzxHKkC9SYMYcYnjg9O6l+oLCCFgEDhiHhCQP
qgx+hEd417JiaNOmgkU52P7eakxUdv/NDJ73RMwBSWJFI1sPY5+t+mLm5XUxRYKdYZWrzhNT1u/4
5d6brr/fE201yns5luojLUa90gBqZ/NMf1EiXjUr6UbsLClTUc4/RotyoFuAnmprtxG3FYxTTkl3
RVu3oeC03xux87c15R2SxgHbkYy731tHW/yCD/tMwkSY+zdRBTTYMeE76INTITQ1X9g6XhQfQ82E
iHOr1aHC5TQFLnr34Sp+PcD/pQN8cVjMapSZAv32VLeVbsXABNH26RMkg8RkvtXPNQOtdcT4yf/9
qsKQ26v85h7wz1BS8hj2HtVWM0rwxQQSfQSMUKlUiQPEpjwJy+5h5dAzS8SdDZCMHdbarEPZ3axC
YpAvB+sBZuXplhtirXDgMp/MWwljV4ir4sM4Q14EqQxOaZQmDM4sSjKbUDYWNbuurIMdIz0Ewo2t
kDj7ol05JXoOrgMeayZixlKPrhqqJDROSwZpn5ITxY3sJDjskGpGcxEVF4KlpKVYJG3+BZuOB0CV
VLpYrmr7ePfqZoTjFJVgvCh/BTVQdcjrplK/DnBAMhH+zZ9z6dSNpZ8Gy5xpNCWaNSYhhBp5//iz
RhKH4xBMjsAcvK0LVl1IxpFUKsJziKI1k9U4cawzZyIHEFpBD5Hsp45z+xwcAPlk5ECznX7PqYNN
YBUJDEPzBmNHJGVGPEdamWTb+IyfEcPwN4TPQglA+kp5Getm/o6bFAltPCqFqfmgf+CwBjOO8GXt
9yk1rbgnorPI6yf86MOWZ3rC7iLRkMbcsTWLLZEqTQONssCBswLgrUPAIPtMr5Uqe1yNkRQyTBg4
ZkQht9Sfb/gQfBnhyCtd49VEeLkyjWdOVnq2ecezD1d+K/Pigph0FiU07Mtw2Y0E3YxYpkvl4wzC
j6muh35R7GexMN4ln5IMdHh7EiuG8Qz73cuh99JUuxQ3YPsu+bMWQF7uqTB6yI/Ia8Lb0RKW5ca2
4FtS1Rk9HzB6WJCBs5w6o60mndftky4JZClGBUBg0hp/sVyvUMghYm4+14mwnLJdEtasMl2DkTlE
5hyckevCr+DzUojw90d4hD5psAX0Jj5wTj4QqBXrYKjfdjx34M7rlo+lir0+mR9Au2z62MQMsSxo
SGf6WDXJh9ViuC6J2BnrHlvTQeh8zDOmM/E4cfBPCaUYShjmkRCCwg6DgBVEzzjIcOw2M6iksDux
KS+bKxAV9sq6bigI0nzk1d1z3Uuc89q9bVsnobxXy5utXF3o863kTMhzFet3PetLGZK9NSMI9dWZ
lhkkf/5IMFdcgGFc4T93O5hXommUeqL1MZ/LyOP4ibH/A+CNFFWQMWhJOFLbhoGcR6APKkk5w9MH
Fj6Or+Paog0MDVcWItA8fNkD2zv9OEual2wVkrchgI8Aqy+cDvqWqn4j8q47D1i/g2NxKStKa8ej
4gryhJ7HGlPbMaLYni9GqPWBluGpdvnBRSWRse6lcLRuiRVb0VM66jqumLLtWXVy5VBrPopZdiVk
chNz7p46BYz5NVHAzLNujBf2+u1U8hdmkxuHbj9Ef5uTaEq10FUtSkkB8J/muFUim/ufh4PycyvF
JDXn1lYycVzvGy/4cBg/bSF9zOYcrCgmWF86zTNh1po7k7hc4Boay9zF4pz38MjI6kWn0LoyTeb0
8dTx/AiIMcKifj5jntI+zCzL3fry0HmohmsKpLwIwD1uuZeNXLXdoBB6pxdchAEm1PenRNEVg9wX
pNzZFpL+NnWsMRNsbOGoyGy3phlOZ3iX9XpEL4aJxqGhEuGSoYbLVHRUm3QK6LKokSdhCMnMfRtM
dF9QyoBOaDoZgW/jHgez0hw96AKhPp6RD7ZlBGhmwQVuDsFeH1yEiDRiYPF2jXf7Azu28L54LBjU
8DMmsyeLtH6Q04w0QP7GY5tEJ5s4tNvMG6KCaPO9GjD1GsuesvNrufBFPpt6sHxLaLlQZwzMd7D9
zu9xgzoRDUkPwS5XcSKkOAn49vc7QxjFTd5+XF/JB227qNnJeSr2KqLKq5uhe0x9woMzuwlAvp41
1KFx2XGkAdK7OsoRyCB8/gab8ByVfSq6GRX0hgpe645p7I8Am2la9+ia5Jh3/Z30C/p8dghv1MyW
BN/wjINhwxPyHrgP10K/wwl0fA0Tl6NryO147WUI9ZKuiD+QhLOj+CIAGJPOt2Pd25uqB2nMAjtF
NNW+fTFZqijv+je2AU3v08+/uYn/W4dE7YBzcu3lT1+l71nA+LCSNE4FjhKlD2mZHZcNa2RXKy7M
Ih0bBqMoXFXaTYPMgq4Ut7hHz/cR0ENXIje7+tAoi/Kv3asJ/P4sPIKXaBEQj0nnQpBL+yhXNuOF
uuNQ0UPbyELhxqK7MNloaBOP3aicVzgoFXe2lRgs5oqNzWla+WzBSCOAeBHGIIekp5DBA4owiFkA
tQbinHFNHcZiuZWirdnuicAcXz3RwvUJljKGx9gmYMdLkPP+DSmhHr7cTwy+zO4XfnBHHnANN8hj
LVUiDq40zAF09cD6C0w09/CKDdrDRS4I8GDtWm6kUDuCQrvaqEBCCAwNwiX53E9ELRGk5BaFdYIH
bylY5qjUrFcTomE3VmU4NemDYYvVtkLb5AzNDkTPJC8qx5ly1CJjRCkeOU/v19YTMhFBCqKdwHCU
HULE8Yozv7MaaAppW65VKP+j/NCk91ZiovOr4NcK2BaTaWoHaaXnR0A0MrInayeaw2yxRwmJBuGV
Lv01tmI/QF0IBEAe6xjv/VwybdXK597QDskbe2Fz6lLrYhqD9BMk3D4I4bBlzxBPZVMXDkmLlWkf
gAeaZ5oVJVrPkdBcbYrKL5GEKpkbZRBcVp+y3PTCX5oBXg46xa/JWy8PhMkw3Lb3Tx0T0vAIp7tc
F+K6AlPRJo3z3jkxJngrFrW6Z8e81E0azxzxVO5h8p8kBPyqESKuK/HbPONSgU1jb8KhlcvFDe5Z
24BdAx9S1y6pjh5+3PuffnrBCF4DjQf5Srdod4Qwuy+ouSYAIR/4IIct6sm+YiSJ0kNZrrwaki9L
b3gjK9N2H3jAjHvuYBOFNii4v6IiIibSur4QHW64l66UD3yIwf/NU/5fdactz100k0w6NIt2ZqFT
mPPsdDdD8BKVWunZxGOtotq63kumWRs/ODEwaIbUWdANsajFlfxlwSD7n/AjvCqm3tW0bkQ59BIG
MSe7nh/n5kox8fVzWRlAlBdHfi6tW8O0JsKxbYIQt1yx9hXEhUfzW+miJGq7hpLIJXU6egtJ9u3k
enXtdQdSWP2sOm+ELyMynL8j7o41OgRi1kfVCCkT6utMjcERcOTE1QGSeMuGx2UgSa6E2pjzILMJ
C7IKy+EIr3PmQ2YM9K9/Px02RadD1UAaDnV4gqHamj7yzbohOYJKQaNv2cr7FFG+Ecm1DVf8jKV6
+1rbHW+UivnNlpskkqL7PNtvc/t5VA+LNfFfCJKsU175IhNm59Qx1oYpDRYOc+JLQ+obTZ1+x5eM
RmzN0jBluIXvmMotH8+ZyDT2NryDuyht9tb7V0Iwa7jCVYjh/YOmqROr1X/9BlxQZFl+M/1t2LKx
081SIEIuhMghLhF8qngbNx0cf7zeSn0imZulL7cvqeLakHTTSNelWn8mMBASTZnEZ+pc1w6YTGcP
Hx9mOXwEUZhmtcp0x0nf/Np+DcFt+9rMgP2wURxHn7fC0SMLCKhj0A+d2Pv6uAywzKxhfViF/fKc
Py3EoSEzsl2phwv+r/MtJpSZbqyhTiB4rsBFGMHMTd+OEF4HIqDYS0mxuPr7SyE9IRCZs8K8xl4P
EBEoxKOszCfd76OhX9E/HPtO3E3WNI8QNEGe2Wp8Dkp/qnz5Iiwq6n+KmYU2Y+tOMFVh7hvprlw3
1BRhsRSK5WKEiyyY7rzYaC99SgdcRhbHBsrL9sbLkVlewEUD07kY2H34GIkbKT+KxEyENk7aDffg
GDlkyVGGbp+03UId9ip1qFHBVLq56d2VY463+yvZSTHUA2BaNCZr0kC6fMveIsQbCNVinE9CIfKS
OKhHe7CCS63rAyk4R4ptdVfT1CH4Aa8cQSnh3RY+pv9FbT7uGzKmOeKqYRBmyQClC94udmN6iK6o
FMiSN+iJbpcn/f5bMRXlYURE8nGGQStduGO5l8M/H0qVb5qedXCLhmq0IirQo//enNF8zGjw+Ep3
YvrGwfY+RqKmAUTlqc553qvj1qLXG3CXFPE0SdOEH6oHeKLXZ9mwYIdkmxzhxu4AvX0e3KxEmIXO
hQEcD2oRJIJumOEFU68YafFzmxe6KSGLKOob8bijzyLrlHRcmy0JcUok1dn/bqc/IUg2/sPz8HN4
HhQ8wKz0TaUNJ0y3vvtUja1z1YOqCAQ7aCAGDJrkKXZLWKk7SnoYuGO77bQbzJlrv9cOLPYizdz5
Uevokw08j6C3P3IcF9U2ogTeTJIRyad+L4VUiWJxE5ju7CflfdILFLgS/sVU8J7eevHAkvFQZADY
92ryZshv30QvPPRxv/LuvAUIxCtAHar+sFI/xH6H5YK4FXyC2teBkoHrEqnKvAvfdY+guuhxCBOw
KyJ3X5Q3IdTaL0jIpVCp+w5zZC8c2yR2hHDjq1I6DVT02MY/3tr4PEBXI2KHWYXYzQEO925NvudX
WzYKeT+fw9Ut+itQhCX6th0ztdPgln4KGHrsuee8N8xBY/q1enOU9N21nSOWf9wQohS0nbnW5ocw
gaEUoH3zCT9Sm3/ZNPdKPnsb1Gb9Hr2puR8oaon0+o7vOm04TROr0fWcokJ/5TlepV6/uc7TZE9o
n1kpPU8I5NfIHEweQxasn0W+PFdlqVxGggBILR4AX1r9EOpDnFy+pUXx5ve5FeyNsHiuRrnLUraU
mGhVzGhEek6SzV6unvXCzbQXoAJB/DlYaWWAaBsGRKhLG+NBQ6zNboIErV6b5JA0lsIud7TdQHXQ
vYR+PXMqbvVQEwtAyFBT7fH8KkjZZY9v2rqbuvuao1ZxPfOz+jdMd3M87sPH6F1gwiSabc3KmSSC
lPcadyyVL4+uztnf2niby1Go388lVwqvhKFhlWv2OhqXKhV8wHHMXpHf0RxpMGGnKqxZ4wlMdWRu
ZsZNPSwBlFgne0yxWSJkFlNhFALn6BW8vp91sM/JCTX5PWQWxXbKbV/Wi30Vy/wxzJSavF8AxgM1
uXQSGiFFYDLkROR6G18fAKwUE+fV8XvelFFkWohk9gZbC0JjX+Bdlajo/eGpgE3Cfb4S9OcNZwd1
MAXTFibqUvF34FIQzcBpccSSzqlqff4JfF3RSzdXPBVaUGRSd4JjQglzt2QwXulMkzq1Mi1tmWY4
SiHVSW63jrYMsqkTorlUXZoqGoPbR9gY25D/0Lic+4mUv+dFjMvY486OHaXguiwXk48BmMpWblEw
eaC8r3UdYguQacUqCQZLLjc+uwWA14fJzKIpwInGYPybZ3YRFZrD0ZBVJ38NO3zUrx3w+ilemvxK
CECGVLx8bmH+AeP/enQBtAqXjG5kRtXicg2L5pSaHetlf4pFNHOaqxPts+YmmUWmnQCca1hUzNPA
Pau3lNRp3+ZNsvkxOs94LNZBgDbu5ZYrM/9cQ2HqV8KVY9kFObZvclgiGs/Fg7gIZ0hUKTlqcM5z
c8lk6Zajlx83tanb8hHJhCSsB2iFvVigouLJBBrqmKlX5N5dMPRsegtRhYKk87XjudTkxksVbaQf
g6hTHD+m8RQAV0Uvl7F/O3rPwAFIZuU0p7h3g+noFU00iAa3GIizzbF9wQGu3fis1pZfrXxmhJjW
NVYy4xuxqbSROpwSxPDnXXsyx0VEMdKBspOqz8eAGPZlGPDj3W50DqNbCTfZ6hZGE8DRwPvP/yMm
QVjpQ+laTgUyohEfcaRye6vAwEATZizYEdgFIwojYT+aeApZkbjI8ypzCYF/DKf2L4Cbw/g78rBc
m3GTq43oEESg+3fqU+Pmhsoa34uoDhtMn/RCAsRC2re1CnCYrY11EdI2SYcjCmkHBT0NKGJGwouw
zhPqdZvKAaVlIMQ5I95kVI2cVfZOBSd15/O+JDqpwMbcYCPvx2cInB38DjLbHVsKOOfYbx14gxIC
5/qR+WYaYlE9p512iK2dWC/0nKmEZULi04Lk/PFhOpCHKqKZgmpwZ7MxByW7uV/Y3qafwUF4unK8
YeYzcUg7wBHdZBercmJNI3k2ooMvk/d5u1L7iFFofwUSo9PlY3iDyqJWnRy8XKctwFo7zys9gP4M
uwsQC0xDKxjSkp0KZMx4VhrC9xErEL2ClCQ8NTH2YuV2A1zntX1qiyP0rMsCu5wiomyk0MWUEXUA
SdAkM0/hA1XB8oHmmzQAswHCxRqfDCN0jCCqHvPRY+657EDzKt+QyYVya0BFA2nRfYaxdY/CjeCd
wmnlnmdkISZSSfMknRvQQFAgHpaJwCMknM34CRJk8ni/lHbQAqSFNJPGjSb1roGI6u3upkpGMzZu
sRNzujg4VYI3o3IuBYUuvXv6RM5u6vCPbqN8eUcaBkgs4n3f4UViPmxz50iLvbDAHpdrMd8MVrpX
oRzfGpTOcdkkPDJ9EDtDPxYEVRhlvdNGrj0cYUTpbooJ23HywF48FolD5BmrstndflAi+Uy41Wig
gx+3O5h2Z3Kx1PCq49KErL784vnjb/+jpw+4WUJs/rNvVEoY2NyOFhlWsQE3Tz2fGLTzHHEZ5QQr
JEmFjzOfAwDJpxgHcoxOUu+tQng3dr6y3RV39+kMQUY7y9DIsWiGelcIIjff48JPvaVa1ttVbaEx
SR/J/LneUsou1soI//n1Ho1klNaSSTAddkaFR8ybGrVHsB41fePNGJKH7AjcWjo9UrNcVjqC6olU
hmUOZ5sKAr2H9sVFxUXt9ob3gRYpM+1xhfowCd/+sk3ExUstKHDsyh6hZ5QkJeqhvfNHAeMelP98
h1YhnwfbvxUsQkKp+My+O6CJi5XT9kUfCKC4pJ1a8Q5f3LZxtqNodGd+owj6ponbvq/4s9Fbcl0H
Shdyc/xmIo6Sx7DuTzqKFYcDXe2T9ghyUp3SDvRDcIzfQNn+x331oiTxODx/RPGkRxo1rx70/6tV
3O0qoVONjnwzl6RHng/wl8K4IXoFpQdTOTR98KF7doKaH5ObGSv4Q6qYQC0YVhlvjVy/ECFuLJ7c
xpKfK+vPcEeNV1o4BZghYY07Bvt3704MowASOWZpvIVTnOaMLVRII89OawjIvjoNMyv/JqXWPxal
AVm5j+N7ltXKziawGbKO4UybZ4CuzW+ekrGLEoefbq6Bzpsh8ldSCdtI7nZFD6pSq5w4DZ0IsZZN
GO9/MmynZD25kD3HFs2KXcMrmLjGUR3ldbmJIBwqB2ZOmjkdCpFcX5aKfDYDU1AYXIUQ3H2U+f2u
Pu7YyM8U4O/UFagengCP0JVNQxkHBsB+KdY4ABFL+DJWhpOc2dJNLTJ//eFMJn3QJNOinhkKwrMU
y5eB8r6Krzw7roRdf7jSlF1hhi5rH2dVDMV7f7Rjvi4D0bd5RR5XmZ1v5L60a76HX/4AmO+NC2cc
69uRAaBjOMGkRwqNUd1HJD9+wXo0xRREthNrv6gzvbzOs+57ePJCG6q4TvVEVaZetQ1cjqCKcidw
MKycbrfmL5i07to817t0xh+ILZPWQkmq3h8bhT+2plQXMzdF6gd+RJlcC5Pkxnn9dT7d1ssOeOlX
yTJLR2A4+5DsVfCm4skQC5NQjFkY8X2k83Z1vAuW/HxZOTvR2OsppwA9rafSeG0lo85t/50ZZuoH
ayYypEldRqMIguoxcQiQsHAABkpWVEEoFu0ybTzt4Q5qfHqFxNchRezbx2yQSoFc5g/MsYJDVMnD
+/LNgM/1y7xOOhWFxcJoyUatbvynDMgm+xo57vJRbTDU7wbU7ON1fXPH5sN4NYY24oLQzJh5Vx9E
aQYWoqOobuz1lGcCrLG3OjI03wW45hhtLUoNx0L5m9Pc4OweyE8e1c2+Aq0UYTERIFu1cn73Krl2
8mDZcVjquyr6e7SgSSlDskaXAOPUVvrmMGTxUPcMlGes+Y0piRkszu8zH5rFgPZt0McHXuHSXNJz
J94hMTOHg1pxuNfUSO43xtlZJL8W9EEtQLod0UDJgFaiLuG8uMItYsSCUo7Ued/OF2RHwVJiRcK7
0bIyhehWYOst5QR3522G1fr0A24J7jdchFb/RfTg48DSBSZBE/iJbkGccvLzHOZAh2ety0d0cTuO
9xFeNrNgpfif+YqzdU9PBPHOUhgl2da27UStDb4sexMDwtIn4/1RdPiO9HOAGErzG9d/xxxiX5X3
WQqHEVgwasoPz2wkCWVCi+iPsoul+hyN/LVGqjkuzeOFwaSlHEU6mxM77ua57PyVLhtA87KljK8Z
gyRUxBE6fDivwmFZIGQFlOPBN6VNYkPUcSfGB970sNQh4xgvTcCD0jH3Jj+JpZJVyn8B7lHJHRGh
sIPCuYNsAbsBwQRk5Y17H4E3p2FQKlI0JNfYDBsvnyR9aBgc0SQ4K9AHbX6d2oa5O2MpfKv/vRZb
ZMLFEad7T949Q3StiT/T+unmvKcD1mLkgTVWc4VKDfF61GietwNGelTC2QhAr/NOwM+R+1d/97po
NLLJm5tm6SrAGQs8pzuTl2wjBDTUIDq3dRc0t9jnsXkMXaq4fPYhU/85wM6gLVPTKGhJoVnceJbB
A8WDNgzvjSAgUD/qchNg2twi/CKNAQg9zswaaJEGlLZdvaQrB4AF9fHyHGwsYMgzwEIU8NAkpqMC
OC5ca00xH9cQisMjzfBMaWNYEB/QJUBZt4UXdrC4udqpXtZ/82h/zxlUGDpN4zVKDFh4lNOAr6wv
AOtv+boM4897abdY4QqH79ixgCzfjrYF5y5fovOX/y+ld/EdkXOS+uJbsCydc428bW27c3K0PaJC
P4i4x/0pICYmpH/OhxK+DQStWOKv1tbiLnR8wrkCBEJkUuxmYSklX3ZS949lRsPO7MDO/sYYj3cr
/oTtSHOFh3W1dNAK/WvOxiF6vc4BCP5tBh3Xx6xY9aQLEA00lTJBwEp18wgrVQLCnDDfIVxtYfZE
Y585Db0f16/NjCF0fh76+HdGh8bmjwmvoYFinTkMM815o4xwByu8t4OhNK1kp/49giDP5wChQdxC
KoQjirzVadQvPWXUhxdCJXq5k04Wt4Qy5Q0AcDATjwzSzvpd7NCz0nCHUcieiyJq+RN7/J/r4hNa
yUhEB9pnAgnskkEvKKloNF7YzTwtxzEHyMkcr1F1m+Z13VpKEX4bOXUsroOJUJK6VUK4gkrjxFgz
E1Sr6BaV4JFiq/A4fDP9AOaEKfXmBYhlQE41kJMR+MYmJbiQURaLiVUQ6VuRbbCo/8icLVXX4nX4
Lo+JeO/E6cAaNmF5A7y0BNiQ0xU4E1c6RQ0hDYRukRUnPnP8BOst/fsJwdpLeoWUbhY3x/3RINOU
cVRjQtdMVuq/XzMdpSX5QL0nOM526/83Tqs2NHh9gMiaf0uckjPFOXYLsMLKD3i/C1tmkccmyniz
38ml7auHueldXm6Xs63UpK0qtL0pg9F+YxQE663CkPIBmkVvoET7035tfymMt0/q4nJnMnwctxZB
11bWYCi+/Mfq9EpqMTaa3HL1ZTjdXDsni62/9PRdTPhLGfzsNDLpFuxhAiNfFPSO02bfV3G03Ulb
HAlfhMrDuvx3dc8vxe+kVyxV3QZQXBpqtPWie3X5V+yWuuPih7UYkdIB0y0ykj9hgKwR3XzCkJLZ
vujzEYinJK+cXq3EgQFsOPaLGHdl5VUTgd09XTzQ08ZSRYAuh1oSkv2JWQnlrc7b/ElsF5dGLZWW
Mf3vy0DTgV7oPXtSz1nzSNGSZEVT0TBpNK0RWPFszGfnP3+1A/WYxyCrAQaSEqJr9Mg2Ju8OHlMw
MjFk7+yypflJqzDm30aLuRp5fJrNJZcFd8J8gaYV68DoK8p/TWYd1C+Endv0uOUZoDecLa6VrK+L
Jp0JdMBm+nxhBbRdDA5Lt15fcs7bm27K6lVEE/WUrxw+FW3NuMDPjHiTWZnk3/0c+GYu+DHXopBH
0IUbK4qBfDSg+3H3+EFbrEIfyKy4QhLOTl+64WOUSuWGJ7wrgMsq8DCuOkDk7RkVejbTmpGPlvNi
9zquGS22uvKapRwLWcrb7+rDYbUFTgeqdcfT6U1yT/UCAkODE/Ya50zCWVC3M4+IOgBQzdGUGgHI
n+iltWF5kCplNnTgsY8eRoJYr9vzJcMTv1GZc1ndTcYjYk5cfhZz6ZwvMJvCKBm6rloR5zlBUKe3
oZzTS0eZsWNb+v8Bt5JtSK6jrOeD/8DpqJuneu1DkSOG9T+CLSd+jPLDT+JOdEow4ubkAzh5w5JU
vO26uaqOMWjc5ya1ekh+XBt385LCSNoqmdVIeZ+UAijOoZYBWl1R1h3PMmBfvmFxzquDtvSaTHUU
4T/YWzCB+DNqPJja6/Ds5oNMvPKW3uMWLeIbLFeD+ug1OOFO45HiLEaFmvOlsOI2hfu23ka/PKft
c1BhepgotRfaQfNL8ww/x8azaEdq2xQTCnjVut1+Fu8RzDdLtYb3ASmEwLDTZTaI7fFlyH5HcFXt
66oS2Tr7/mf94dUX8vKjivN4PaxQRwhccIZFs2LKB3SYs/iPmZ2OR7YZ0sdGcRgmuweNKHy5GxfC
R3am7SiGU92/yqiIrEXbRyjDCRsgIIH2PZuZkrNXqb1Yhgo2M3ZG6e3Zy8UUQiYtq5rsCvP6ViY2
qW9tKs4Ryo22wcqtX9KO7YpVGJAiePR7GR6ZGV1ZguPxo8dGGtJ7CJOBEjtZK/OhV50PsdRb58W0
ykUAmp9QzeTDMU7F+AWR9O0t8v+TeY9C1wzg0PtORRfl/nMMTs70Jaw7pxbT8CZBlWTLLOpdmGDm
d4RNo0USsFSR/scNHnEqgxbLfvuYDCaGwJRV3XBzucFJ218pAVHQiZUV9mOCNCy8vqe9ntNtkgQ1
+FX/B6y/VaR/GAlQT2fOII0mUcPFAxbOSh5vtauaHUaBnzkC6J5AnrEcTW7xHK3ZDHVygFNH9Avr
ySwf1McDltXEB0j14myYpXE31IjTyFNr8Su8bRIxCxdxUzqjh63ns7nrVc/2nBNMr2Zt4gIP29hj
GxpF3uje2TV6r0oYrfk8SYQvw5oylRntLKGsA5LWC/oTZ7ZKGFtsnewNcyNui7hQDLcg9R7v3OFR
IGdNqTNHhLD3zMJq8ZgzvdOD2j861szaPh8PYxBZ7SWdACxs1lA5i95l5ZeVCn81hQUhpdUFP0KT
vkv/Fg6EmwikP4rfdsLPt4Ma3cwZFFgJ3vfOg4CIUBgwwJMV/jwGBHB/PiIm+ceWXSXd+Dqa+wDO
KwRw0SnWRtDqtfCsiRkrjehUPupWrf1RWJ4T+sllARknq43HxoSlUc8eyrscSmUndMSlKqYaNtmk
jQJoZ4foxx+lgzhfwGuGAxqZm9KCDOqLwk9dQTsLwkcVikl/CLOfz+KO4uHNUZhLRtJpDSJInlqq
MFd5oJVOn2xv5AIWU2I8iJQ/9cNgJcD5swSQP6GbhAm7kjBQgEHYz2F6iKl9EcYD400P3qGQaS7a
NVWGOBqNIjpa1exjQwdCoLwFQTi9lPhebJ878DI9pQh31GBcbiHJYukMSDm57EaQDjWH0M7j6Ack
7M4SWUb8KSN09ZaD2SKMZ0PVLdvepuEbwzBYZM2jdyDiuH6xUrrbQwwLCsTbNWQ3MuJYOqzbUIG4
ziLhfgOUCmut5X3Z+tr+YuzHVFRmV6BcJ/6W/Es3oU52Np5UCAfXnQbJQwoAc4z3T7MoD86AScBq
ual9WuGdFiPLg8Em0SoLlRZX2JhX1uBSxND3rncjOjk9ubWbaGUy2n031Ga01a6Gyp/vhA7Wys55
TNi0AiUbvzOpzUR3aCsvYQvkywhJg03vrNEHiK45oEcJ1jDm+u1vYRw14u6WKel4ULKsFLXkAv3B
mfgVLhOIxNWw1ZoIKJXH0pIzyekYDfVn2jI/apiAJPWxYUG+R9eevcrZZttGNuvDaYFMUE6zk5fa
HkBgT1mBEHLauOcWbzKxyjpqKn4HRpk4y2KuBSFN7uMUgEtZJGIgEIvQ3GSmYRuIfQFngi4wxEp1
Sr4+Td8+0GLLNSpJeBjMS/70GPXcBPLZgSMJIgvibohIIdW6h9I5lTpSaXJ6tmLp8eLLVMTSgL6E
DyEcJK3TApIUjjwS21C/b+6WpSnIGvTLPUksTVhgXeL9MHuEUeycGE2E0emMe1xIHA7uWkVDaIkS
GVLi42ztL6N0OSvHcxyK4a1ET+Ay7PSkhCNvpB3F1TTTElJi3MxV1nDnkO3ikCl3cVK9bUhaSubN
d4BOd3x5dQ8/Gv8bYFix6dWQmH2w9771gy6kGHTYv42ETz+opi/rKiEQEQfk7GpDN/4YxcBsKkK+
hNRQ83f6OuaXygoago8wnN9qqxJ/lkHn/3VsJOldrWVmN2Ms3QKHy59vmtomKtla/qRVTQncsvK9
K6B4Umf0nmH2cA5hhzcYZ+bX8w9uah4PGZ+H+fRNOT7iSy1Wm9+b0+q0HvTkB4DrJIXvbfCY4Nbw
kNB2etu2G+nH22cx3kca0HRKJRCN3wmxd5mGDbApBdheFmnfkEDRLgme2qb3iPeagUdc2gQ68Jje
J2DsLD/rLBC/4sj4pjO5jThcmj679PcGC8Xl5SCkupffy5fOinFOxnANW8MLn1toC/p6ghqJo/sK
J/+Jp0Z3P5daT0Pvq9Rd8MSXFq8RgcM4BZYBzcl67JUAW4KVTBNQTv39dWIhWva9RvKINK4f2skD
PEX2/nSQNqAPh3PcNX0IBl4YnN0COnub9rjYLrcc1yQSxxXNjUw3tSkW5GyipJsg07E9QhUmCWvp
QI0ofIwtL2mi25KECjhoVEsil27MosNJpF6TziiO8XzwbUub61kU+VgTx5lL3ajAXjY1fPNYJ1z7
F7uTK5/j/6uDtADfXekZbjw5d9Ujd9PKttyaUxtJekBRMroQ1RjvpL6tpS0xVmaZRibZx5eNXQb5
l9YPZj8VAVKLeSHIsfY55FK5/Pg+ozpPV/s++OgqCTIM12nnXljScpjvvHsd0zGTK4Fkgg6IYUSR
dzWdEww0YdxMkY291qcuu2rK9wmo4CJEW4h6MTKMZB9ps0cVg8qTkI1bQTXgCvn84UUs0JXY1HAD
1WWsNEbSTiJq2vDxtLqPilkPVjx4TDKZ0yEhmz+OiuTbT571+Hw4AgDZKWYK4y5F6bYghaS7vxiC
mC1bUMyKwNbc+0RdMqMsBGiB5/AxuQ41g8OW+ZO0/8mYvAhGlPQ6Xf15iUulpNA/QRNdtCz+HoyN
ZX1HHeeTqyw3yZgTdaAQug8us2NGU9Ti9rYE6t+Q2UaMsthaAD2CpOlKoQ6dDP4j2IBpWGwx8HMf
75MvCXNYav+8sAFX6+/spme0lWMxLTnZU1lbNYDiGGHSfUR11E0J/5PRbRsIQEGpKItecq8OKm6E
ZLTY5iXwmo1vSXWYjxuN9HxHJk7wn8vrfcXIxeCw+1FZOS7/QMm5Vb6dESqvzVz8iJjuIh9Zg2Dx
HDuHj/xBjX+sqbV59HIvXQDwbk3NbDHubNohDWQO+LsZmi+1M9R/z3sB4KahmsT67oKcCporxM+a
SVc8SMU2+hVSrcqR/02V3j5M4UYcpzzCuFEYj84yYCbuVU+QthK5YTePrLTBT7RMJmHTCZhH2IhG
E57QFdaR0HBoe2lJeA2FN0ZzT/zXT3/YvPnjG/zr4Ro4y0LOzK0PmhWUbokLW7KKvkimiSdZi8Nl
UC9y8r3m1Esm2SF2m3QyWh5qaTdwhPh1/lPCu6K2hVFBXxq02v06hEiKioBUUsd/LYw+nDzzhtyD
tEp6Vu+HwBmZ4Zwt9TXoSI89r6ceT+J7nmS4XgrlHDqalxruWeq3lj1T7Go3lX2e/g6q9Eug+8Fw
4H0nIEdcUGtqboiXJQmh9iTh667RMpw8xvQ4Qug9sleHshXDCRNPxOIgVCnKPRmkc+eZKclIzRW+
84GLpYE88aav1p/Pg1zIoi74s3dSLubi4vVXEWYk5JSghn1JZbEV4GjmLZUURp3PJaOXdVL6sioV
fFxCqF5tBCC1l4yxKFWAxsfowiDIbA2vfYbV8bRFK6YImVG+iOqNTDJTQZooAtA/JnEA9Naik1+L
2KrdAvXOxjdjw2+Irx8GRU4Wo9FWxNQVuxhpEgeZ0Kx+YsEcEFXD085iJ4fpeTSLHZbKnH45pOou
n0deSopBMYdkCYdycLVaVbPmC3wIEIN9yePT2ZiDtdY0wlJaFW1kenrE8L/xYeBbEaJtPHytVtMH
cL1fOCPayIWOJ+CNbXc2s+gViF53OrbyPdnlVLS0GxyWpRuQClSASHHzgJSGPn73IYY9fnzgrasa
BTJzEI1/tN+MTq2z77yt3cg5xZbSaz6jTsrrw8eIp2Ud9oZ/Z+X1p+mjW3NG9XWXGMvXFgez9Vvs
kIz0LhRLAxrhlMYXoqmdwKcax5z6TPknIOQouiLkjmrXbyOF0c3tGX4jJxa1pshL5MoNNIZGS8hX
2TToiLeUHpTvFKr3Qdv75OxYnF9bsc+fWEJcr3CAmWy0XQ4vS4xRif4Nwjkd+p1BwBtI81w4Rd3k
XnRtlOndo9Ri9TW4VUclvC3xv0tvbFOALicDV7/IpLO0XCtXMIaNaN+oNP9ZRgCIYcHdlN5PtKRx
GNf8+f7EAe2lXL0QJrFLAdo27pm95v9TmUTbhn2uRmLx1JtK6aeJQJTPem+yVs6CqiiiH6q4Fa2E
CKXqMpkc7LMRdGFAktYJUeORgh4k3S1nEG+ann7Jw1nXtfMAicyyC3IfrE32AQrDjrUsXsp93Wur
A5E/Tr7PR8FXwsL3PeP++q86KWGeVOdgMIBAN0lC5ZJUnd5FW1q+zar3vfA+PRdujlAYBLiQKPkh
WQDoJK/VqPG9S4sHVt20Do2siIGrLNOJ4DAv8plTMufRjduORLolykHR3wZAvrUdjMsh5efV/0ai
mgMYKhWv56jESE1eUc+C2yjilPIKukl5Qqhz6auQz0ukABOITSpfVLGLLVYoWPxwRwUbJFDUgsZB
8CfCCLDzym0uIfjUv+4OCKLfgjnjLz5QjaNIxwm6g1lhvXn9qrOylyvHBDqWz2QloZkQRc8nqelC
R/vnRbKyu/GNtctE+S2Oqn9bIqkbNmt5lUzq/kr8Cclcl4jdB5Ne4da1PW9AkoQQmOlj7OTO/MAI
ZWAVpjgjafKU7XoQjQNhUwZtm7IBGIcdqgZeXSklbvzIec3enBoQQ2giYebYeERVjaWBT+xRFPJt
nYqJwiHx2m9kYhiZ8vA8v6vdThDjarPB5aXC5vYTrZMUHKSvMmG0EpeBumETyccoVGOwoBgoerib
SouQcUEzanLHSUoihjiAIn+XMmKLlyeEFBjod5O5/reTQDA1M8yX1kQ6E0VQaeoMCXN/gf1uqeqJ
9K+O6lpvOurm3igMH4lfn5eYHdvlMgtKItsBCUTwBq3WNi8cNr4yTRM0hd6gNM1/IaJCtafGK8wn
PRycPoG4UWLeF2UTK+TPR6m78cj9l7SGmg2XTHgo3iOvbGvqaKUSLSy4qjK2tcblZaSD9T9h9Hxy
I1UegTSRVoc+7kSHzn9auNBMMd5P7eEpTbZYxPLJPDaBh9WUAuVPLiirarX0MRocBj7NUmt8+ZZ4
q3k3P+T39KoOiAxoRIbG2JhsL97yrUkY1x9VAPNFmqDMHjnFfEz/pMPsnBD6caTcz2wv52uuH3zl
GcLi/MjMFCCQ/gpK88YeKgUxX4on8jWsmLL0uSRYHyXZAgly9SXICx1PvtNSEIMByBWknvQi+uSL
NHjJZbG+s3Hmyw+31PxFWCwyKXDria4IU06lOVhCT1hcTE8fRFkC1mFN46MEVAHlS7n5lnScv41b
qb/3cfPs34SaqrLumgsZQkvvTzR87gaUBGkJv3d1JwGRCNAOfvT9WaaoPnenc+WXUtE0Ktw/Gs5T
pUEmmqYzNziPD5cpOr7V9vloIKBfd2daXUSHON0kW+9Untngr3w/79tBreyzwSgnAob92zO5j3Pv
CSwBXKqBXiIGkE2QwGOpK9DdTdKhGUUuzC/K5prNP4nh5avSZvu0jH/bdR0EM7q17RrhxTECFDbZ
edAk3GcQazOSTMW6Ed11pTDVwMU9Oxmmi7flyJPkAaOZqPlAdE+tdqF+fgLKW/KHhX8PfCn2wMUd
dYLlX6j5V0s965/94bwSqiN9ZJOJ75Ojf6AhskxqQCWraPAU3veI+Hj3CGHciTtlSmX+lLL1yk3/
ScTfMF7Kvwf4bL8sXIl7viRg+J82pfUlBT5MN5UOmqyqFJJO2xoejYrxwvLj+hfw8Gs2/S7Y0gbR
UliJ4gUvG/uH6ECdCSHsjhRLbMgpibkwKoWlbaGoCiZoFLmKa2jdDnV+NvbA1uiH+CwH1LoRYzpB
lJir3qx1ORSaJULXvQ0tyUAMu3b+1trKXHNc01jtTw65yGiPQWHGUh310rMrVAXqmJa6TTW7rJxm
7tpGnnGJWh+CWIifsn7bOWYLNis3096RI6eddH2ibUpe+2HcPxRJh07UGW41vaSQn9hMdkfgSabX
S7WldUAtVUMsyMwc6NwW2TzHErJCK89Z4GYmxi6o6Bvj5/3G66IUH8Qoj7KkQiODpAxXyfpSQm/o
RFs5am5V+OcF9JQVz5Nv/z/V4FknEUwYmGumsk15aSsZa4rqt0mWeeHnoy0xU3IwwSSVjjTb8nHv
xfG6SuaaGmgdIeb19/r8uM72zHxfj3+FQiMXuJIMCQuitj2iAB86qxrD7/Z08d/itVk/R+nWP/Z5
YBwK31jaJPAG+SjKNhbr6T9m1BZzYlmkWWDdXUGPNoY4DtJH/i1/yNpSb8MvYhP3jZhcoGKPcJ++
cSia+WyyRz5pthD+szx0349iYlFI8lVYGyZpTqdbOHwkFVc0STUz+bcqaKCym9mP8nZFvlojVRHk
MxUE6owlEDHnMJYBjrVxHWOYY1lYkmV7pxAWPGIQgyW6YrHCg+VuiOJueRiTxL+8Q9q04GZbIXvm
cshya3bQK7uO8jpg0Tm54nBH7Gvx3iP/G9GcaiyHQzpI3yoH88fflBWBAMCMGNcZNmQGguOmULYX
6pDSC5lqTt4DaK0KQOFIAIj/jUh5Qw7nFl+ZiRVw4O9UEoHeQ2SQIlu1ZjyzUoKQWgneIUDpefn3
/Eoe0rzso+42OBjG9U3An+OIr9cXR07gwZO9vpjjwCuAoQIXxZ9E4pXjLZtU7uKSN9clAq6MCov3
BntPPyzKz/trwXC8tgnM0JaMDD6kAhbDHiuDKI+ZgsYJRZ1JTDmxKOJ7KnCngI1CE6U+8k6yKvKZ
vUjxxO+CaNSL1gQD/ImG5/yyuQceCaX66XgNgyOdSQX9CmG7YOW0oeoo3/GwwJb2CiYLxAOz8eUw
bTVbbF4tEif0ayApZg80zjnSUu21GXyavefxjXFOlwv/2HsMWtoGANNcq9VNXa6z+X+kgX6/L4j6
kIQ3S8AVfUnyO32dqb64VBHEX/MYHEFfdPvQaSSXntJu5SmSAqmZjNDlQoGE012DNldxFQ83wfMz
aWdLu7HyFwEWvLwtb+TI4TqC2Lw7vcr+ZxuqlWYhdXZqiTpKw/IppaHnaojntEnlbfIgTfOCInaU
BPe723qTh2NPUUScA9D8ECXb9KIaaLMrWz9c8Bg+D1hAU+kJUDAX3N36l9CY/kXnerLWUyVDLXxv
HI2SoDpPFeGvWYYtvPyeXFdOkk4OTu193wKgvm3Ku+tMQ6aoPczwHXcr91uLrgtcBYAOcBbeDAd5
85T+P0UuUUChzTsYVSjqc5Drc3o/rgIqclXwLGrD2M2oeQsMBfopZFSw6U81D1n2/Ts6mF1rxNk4
gl2hQgcrd7+l0GZp87NhJ949SUEGpAcIJ7NOmwnkyabp1iG3P1I6C9Yq1fLbXpEJxpd2t7rzNQxS
RJ8+yA/zjCIaRkYJYQ3MRIhhJd2UVLBCqowM23jbBkI6J+txcptuSBavJ/EnegmM/Xbwm36quvAf
zTag48MxvYCawAXVw7V3k7pgKPsdWmmYGGeVc0gi5F/hXFDLYUv+/fn/dv7QWUBMvMlymUHlaYlV
F9LrRIgN2frBbQJVEVMeCwVdyIETNZvkZH6p1PoFDLTKQuZm7yDopL0xFClNPwT666Lz7doN1TaL
HG/VSYR09kdADdCJaW7OMEjsaIzAYdUlHy0XU9Iz1MTkjVPt+IC7Q9qBvCfPlQrir9PL3MnpMcZs
bT8UHCwL8b8CXzIZHW1GwrW9sCg/mt+KkNs4ch34qKIu3TZ0KwUm7K3fJN8bCm28O81gD3tjjZ4t
yisw1trnGRTSLpwXlZTu5dheW90UtI4zFX0hCD5j9ZLvZslPhHtth6PEzOyQnj2qfMaCi1lmWj3F
TnVwH65Rpb4682NdCRNcSMXQeAH3QMXBQInkgAD6rVe0OTnzYP4xhqmAcFBFIRz6Dxf2QYTBZ3vx
kliKMtcdNnh/sQrVHodtPJLn7n1NhvgA/Tfd4nFPz3t2peatGaA3RXYEQ6OSWilCELA6PratE6Vq
aJ+t2E1S6P0SMvNp/NKRMzWZVs0gFsEcDZ/hZ1kc8S8UMarnobKsA3U0Dig+oCwuQ/73bLoTi+jB
PTbaoA1+jdcQ4mRkusTZ4GVmoM6KMn5h5Hv0my1+yNBUezekmZhQUZp/kFRge2gkb8j/WzlYEeBE
xPQc5dk7da429E+nnF052nN4ZC5iIxdfosnCYpsoafOEftmtY+wDHqtcC966pFMzc0MdHQH8Ydwg
ndjPTmzN29nmxl82zSuhjvzPr9fFYpa5bV97gdmqem5xmEV5NAwIYVhzGUvLmlGTmgJPFylHA7Vt
wVy7honH+4H8oHfL0LZFoaS+XrMYD+zhaZkAL+iYLU1igu5Ql2McgJL83PRinIkiP/zpsHL2bpmq
AAGDQ57QDVznizyy1Wt/QGVsJCkQTd38Zja6ufTGgH/VeWpTXayqzaxdysvXazdWSV+Zon+idmx1
DY+fUasZRwYniUONZSZnCuCo7iI/iouomn/AdaIi5sgrnxpy1SR65LiydLLohKEphD6k4uitdPBd
ziaST9I1v6dPo5QPHRAIfFvZ3vIXD4g7NFPGVepSiM3SvbxbeSz/cgz+24wzdSE2frhVDtt+BUJL
Wf9AgK3uGuhMPNRVxijlBE3FxmPHpIB+Nw92alpEs4Zm0nc+RZIi7ZiXayqcZW8GWeF7fFsXoP11
5nyY+93EaUZNwI3atZgPpaI7627V9Bbaon0YkbY0i1cSXBf1pTyA54Oy3OCcG5x+qKOi1elzooZG
cBAuED0rzZ+B5gJM7xBMILOEL+c7txnKTv/rInNM1kx7c5AQZQCR82gx3uAl9c30rh7QlVWXs7uT
E2Ri0wo5ZVmHYzhBnZVtr2jMBqYVy5dOBgquPtQwbbpn9zRaf2uUoYci5UWXx9ChShpcszgl3MlO
a8RDWIcXDQiIU7gHsrD8aIKk/7h+hpunyBkZcZ9KEFqlOcFcQkeIVZnEbN0V4JJsSoqzRQZBnEO7
IHia5W4bkoaC/3dNrd9l8TK/m/gqgOudwjX/IK0KFj79oJpRnvoCYWtbNWw1uTQbfUFNmuu6gcJo
MYPPg1fkdG5k4qt40jkgbuCmMZiH3audf7wMmbQ2qBc60nSKzTqfdiROQfyV6l6oXkYYODvJ44NZ
z99ie8ljQSP9xm9EJLw6Qmnsu6cnGcuLILyJP8UNiLGw8zurl7xR12fu1zDbI9Ki8TYRXC/OM5Yy
omYiP2HXj38eyVqp+RsN5plfsQLI0W/01Xf7BfjcZzjFzHoxqTiNerTwwmA71i29fT4gI7newmyF
H5DPWW9/Zg4wBSJrqZ3Y0PLG7EFIfsU7ksLz31tN+fdjaQUdOEPFA03fjeTDRVcgOtGnbgXtNEYU
Xjj1Omj2xgHatRTjq0TdYPDlEb51fMXYNI+3XmyoEajsQJShcR+hl8o9WdLr1oC2ygjrGKxcK+Pp
fDIP0O+4fSEn/aqwBqsONaakdU1SBP6yN61RoZ39WsL0gvhcM1ccfc1aW6i1CJBkbRyVeAM6cPIR
BhHGjAaepWRytxw60IygaGr6Pz+Gej+h2IDJ9wUmp1MAUxaVEXmy8xTj0DFCOmLGeuclZ+x9N9ld
Y0kyVg4dOPwK1bWqhVYRb9uqZy4gyib6RNwztwd3yUKx1NMXd1aTPUjBK+3ypbeQV3e9SO6Ox1k0
U/bVIPYmXCLUSAwKe5L8qlpI6FRKvnrZD09DbM163q6Tumlp+ITyCgOxLtpRONGpnQAz0oZEvop9
HRO6/FBqioV1N8AelDdvy2ShUjtWtei4FcSxIQIJYIn/AKGwYBuWqeOtBWbSIQRhR64pWK0DqdDm
A+oWtJKOn8YYbeq9nJAdsb6GRcYB/KTGt88wIG9wIpwicBW6Qp3wUyEQs8+jBZ1V9rUr6azJAeDl
9diTBwyrz6iMkMBrhIl29PuWl+xr9wgeIuiygnVpwTaKqI8b/e9qigR5VsOE5yzW+hkx0qdA7KSi
CPlPZPBH9AcZhfu0i98PhETeht9oR53TZTFaBzNL8EUdNunkDLgo4ErJvF5frgj+xXnI0hfvujBL
IO7bnDrNxvlwlfQlwuiCx2fwlEkECezym1hh4p/8y43eT3jreYz8ydzvDNVyEk+UEnx9RrpEEBTW
EAO/p8BWKe0vGsTqBNUVh3oXqTLjiZ/1q6dpcDUKWMkopOpupB40FlP5TaMzNvt781NChHqcMfLS
tLI0r3OxhSHPl7MCZ4Bi9y0rbH8Q32tpAjhQn8UfUHg8aMs1gycy3gT/iAFkIShZ4YHSY3V9FUPP
hGDJCrff9wzIlxT/4St0Lc4N9wfA0JYo5TZ/xR2g+iEbYnel8SY7Ztk3naG5IC/xBRF0iC/d5nU/
Ws328AuINVvw2RYNZzK+YhpQjMajODWA6VBpbHN2zFOni26f04PacncEzaIh5CEpywcB4flGr+Bh
8YXt+U9IQ6WVCxpYIzMcGYijHeSYVOIKqeBjKYa6/LY8HQrniOYNMNNrw7MUYf2Z74sVo+OdRag0
fSnrgU+T2mHRHDRVWyI5gAnYByuzXwpCeo5ShmglzV8jnfvpBZDw6DAYkKdFUR/cAE5Qgm0s6Jbw
AkpNH6SmpR1rnylSYR3gOUYhyTfC2PX+h9A5uEk3yD8AXQ46QEtAzz8xSNwcM35+bfpeDHArZZQR
qlQ0CWfEXXXIw/PtriZO0cyF63/seKO+06rx1kWeb22Pft965l/+4GEL8O/IEdyin00EC2lyhj/0
dXQX3EAm+rZ0yFgg8vdTM6E+9Rih5MEeYnCP6tjtWFqUnD+ofvVJ7GCidOYt6UCxWj1CaiLin0eW
iETjdlDpxlhEsZhoKhFBVeFvJS91rW8SqVhOOYheto/WDjRx69pfpknXe56EyU7U9KdvoVp9xIZi
P/SVi4/t6EJo2wbV18dGgjZNmAMqv8eN3JKwwshQMD+VxDjuI/syP4hE3aI13FoDgIqinCD4rPH9
NrjyAqSZsh3FWGLkDLDGMlVMhgckshFGdwYbkYSESUj6+d1L6KNsjYKRKSG1AGgEruqcqJJVK3fm
WqVck2uX8A2SiVvlzU2ApDTBtSS7QwPHRsc/96UGOjQwi/jIuzIMyQzSECIxylTw2QfOPdUSGoBM
UkoKvJzowfkez/g5VsMXD4gNsEbXIjZAEJEjo6hbe0MPTQPnxy0u3j+1Dm1pihAFZ0mMM5oJtd4s
0KFd8ohSrpLneX6s1XrHZOrtEoq9+eiOonXq5pOxT1uLMtyl1eIbPzWK6bJznjLNSjMd0IqfecBi
hTs5hHgmhpm/LZtIVEnerdRobtzmPvd5M3uGjmdsRqYcBpCN+HZCotrnXuTgNEPYpaJgCYm19adg
EsKihM8rBJvCKa/6rCAzvqpVEiCgBz71shEwY8L9GpUcIUlmlgK2xFpCKBHcEYokhSvOdKGFF7ec
IQCEfUtl82g4to/QrWXN2jO3E9/deLQfdLh28Dd2hSYST+knsYF+LAzLj5MlJkYdBudOIhNfRL86
DkFSQ+wbesTIRz+uZfi2/emKy2WYMWJinobnDTPV4BLFSUTahuPKdMNUF1K7LAFbw3unoBBxCETg
2rYmcr0V/ws0/pQOM1ay9GRMxz/wJtctxwhen/97CPYfcRw7LFnEwrM7VVu/vUyEQ9BssIvjvrwR
pFsUBT+cw5dyZ/dvCal6VZyR2QzH1vbm0fAaEC3uJzBpFpN2JRnTDmxpoZPW6f9LpXFrctHx0CyO
Tv8WUU5sqj+YOj5hLVSBoz+03Xr/5Kk7+DQf6rvyh4dhljjJUi7/tOcgRFDYzhrz3yNvp1QxWlKe
QzcdOhirHpGJjeEUiSsZJoO39wp4CelUgm1H61yKhgR4FbQ2FKpzrjveEEETqT7xkuagZwCua+8Z
PR6u9DOpCZ5CD4yOVF6BSoRiRwSSHhmu1IzLxxvU2mUelxOxiWsoPnNXmf3mF0Ab8jW0EDGea5v7
15eRq5G3AtVfGfeTQpt3HC2u6yK4dLVQebC4HoHuehjb96B9kPw4ZpedidMn+XZwBDheaEFCrZaT
+udzqKx7ysyUoAODE9abSsm9afphtE3puWRqUGH5ecB5my9lVYx0sVvw4ycyoMXLrERP0mtPNLaS
1TJphCrSbvZIpahc18idw0+VaqhOeCns8XheXrEvm4GniSd9g8LyBCSFVaApTE/uXJz0OPVLNw1B
rNEWdjqmzbLeDVFY9PbmOxDN2qEjfo2YYkWHKmxEdU/OBta4Qd/20ElLKx9cgVOujMJcseARGpq9
4wknDy+LKcnInPCLoiiXgbJXv/wBdsSMzuI2Ahdo7YwMdcgmbC+GBm08ZZxEJFmDYmLT8p21829G
yP6CP0//QnGd2GgnlO3TXP1wvJCowgXBtiZyp5w5YdCRDr3+Zn/nM1wWh6e6Ktgv9FOKbZ4uH0ks
oe9jaxBA3Towng4YS/MHg8hYr5e7WV0DB/gvag2M2mabFQmHwVu+Qqk+X9acIiurlOHQl1zPyMpT
ylXdJ0D/lGEvQbtfZv/aw9QOs8AEYdzq7H5c8uQUzhLsYCU1KP2Q68Xpt5Ypp0tM1m6skI379wd6
087qfaiWfUnvgtf0XD52gj02GLgyBwDvk0zqHYXHo8mOvAo2xLvpYQ6AoXeHYDSyYON5PH0EV6Rb
Dutfm65aGSyFYgqnXZAbg87awyanGcs8tnTftHa6M+BAKZdhmiFzqfK5teFd15B5WZ3RncCsnt7k
BW4pBazKe6ZtRa4yMYXtDCSi0M1ETD3lW0xqRrBiYU4muN+xEupNzldNGeybXghfYXEixafXqbXg
d3CS/ImJuscP7bL95zRxFCZ1HQOFdp3lngtzeDnOjpbNwIpQ2O8yM7wAad803znml65cSWEq6FDx
dnM6zHfkP0ZEZZPl55dGRzWKxZwVRJtgC527vNr9C1zYWzMdvRqgXse9EFbYKBA1V9PwPTaXUUjk
2LkM5Z/lkOnsE7mpbf/h3JCizQ8cK3jKHlnloRvKf24GT4cP1l5jGF7mWqUpFzVO47OtgkTQRrVN
LXHIhU6JRvJ73n3It2AHJ8uRWOVU7ioxvIJtbs9A9TTOzS+NK9e4s2LxYJadeF4+UzKRssikC/gu
Z28zaLczy99IFW1xV7MRsRUzPSvA7rZJBJPDq3vgS713ZN4O3ZIWBMdT+Y3PY/TW54TpA15eJ7o+
0guYSdsMK/KeTKVQ0SO09XDZp6ExmnV7/CvL3jL5otAhg6/GGzFJtjeD5Q9C/uJSKtE+dc79x9Cx
tV5+GBlmFkBCqrWCNveUaKXrordi2nP0k+m2kEMUG2UFB/njgYv1T6NnS+CAJcCK20TrjRM6cR8X
IVUY4pTtuu+KyvkKVh2ogdAgCyngIfl11F5kfHmZ8513/KGA06QJictz6v/0LsBJR3hDvXejiRd9
TuJqNNFqMtwp168GLTdFwnAyFVZtU/V3zwCDUusHTM67KfFBMztf3ACZSQNwZO5CermcWBD9ObgN
2VZfWj5/3LxL3VF2i17lSsQSLiq5bV+m77FpEo1vouHYGJi7ZeVmjb2pzhR7F366lHCtHxed3veC
1asoq+R4Ud8VABynq82k3CWgWX/sdnJ4kTFMzJKapvWBvo2g2lbvLQLOEKZX0/aTz5EbePX/OKTx
mpoC6Tib871Ie0f9cU4aCtkkvo8fS2BZHFwYCIKmZYnkGSgKy041zpxkUSsbHnQrqQEqnBiMFMm5
lSVg9RS61ZCSpLbZ+AvyT+Tk+KexwOlZzmMgIcAxa0yX2xUkKRzCtpEaK4GpCMPwZCD4Ixq6/zBe
Wz7w8ZFbHxtRHFjUvUrQwapPGU7tyJJQHPrw4N401zwg1g6TaOt6yBaDUSH4vb1jc21TPX6b2q10
xFfJByFT0DK09kDdn0Ubs0qpN5vrtILPlbgL7fbvD5t4Ev7yWCK9QxZDxrcHos3v8eUXG4lzyp/b
0z2xqRA8VhD9VmPHOJ/r757bRJ1PKeQ1MssZAmwRNramcPlqSnjvbTyniTAqddKakuPML3L5L7Wd
8dip+vVikPgQWeCgzyeA7tnNhcnIdqxyZGP02KhArxsKmV4HXrWHF/lwBdHDhG/Y8C+4VfWHq9bK
RSDO5uk20wiUTIq4Tr5xandTDfYZT3qoe6CZz7CohNEI1g3e26b3dFJQtL7RvKEnErMmVc0xo/G6
tFeCCWF+sgp0X0QROQ5gi0E7GGMqrDjGokShYR4p1FeEjy0kzkpWClLGyR+TkUFr3U2SA4vLiFuk
AuaEeM4o1uUZg4/ae/eeiTqu9SqGMYk3XddmCuL8VyBWCu+wprAFRibjOQF8/RtBWKcIciWD3eY/
qDQgZwa7EEgVKRnaQOFgx0QdN0GOqKTjqkfJ3LBoqYPd2tHeJprYL4WOVN0h4B+srY9bzDt3L0mW
f2woX33F4WPdag1qZuG3yOdp9YetQIqUmPZ4lJ4tDP0MbSpqrh79y40VNeYScQZNer77g/Rc+NsX
5sy+O3XSbwWnC3FaukDhA3fdcqbvUr7IVpWHfGjKgCCIWUSSG56EkQ3oq51LBiFjNKRFlhNzdqea
h+rSlXCMt48VyoohT1eMeazKPyU56jIg+ONd4gdso2szg4lfBshlkvLx1pH8Bi05ObLSDzCGYa7b
Ore+1b7h9dsXVbB5v+QhtoCzpPcMxulqWR4sFI9q0G7WUEt4onpr7VBYjBBJcZIHFUm1/CIQobGH
sLBHhqtXfegTbuoKCC2i6JGTk9IW1GZlch5KRn1U6/7A4H7/VZNVxlUIu7d0ntY/XyWrj5Yr4oA4
73OOV3f5wDR0aN3wteXQMTyAn7djqFfA08Yn1x8d6tAodrroHbaUtDcu3GlXb2s49KTxgpdaRLPc
p5JznsTG4pdXz8jxPgG+mu25bYt3AVbdXoSCfkos0BrylRMKMqBRZ3ocF9ZfGbZxGKjRpXq5odFv
46oLxNnSuBU4N7XTMp9Ca1VcPp4zHH0SVIwIlG3+jThm2tEYdLMTZx/4A7fWHrsvRpL0NxEMRzmK
gxR1tz7H3HVYyJACj5oCpZe+xvk4uDWuLai61WR9DAAcXt7t6BZ7LL/XA2sTUZKShffcNi9EbSiv
8L1q+/gIQqZaiqWvEbrq2bXXDoCjwPzvU/5S6wVttJflBKQA7E5Ip7Ltv5/mEBbkZA/5JIoPaWsT
uKthz0oEaZtxZ7ANVHHJ1BJpfVYU/2HzcYtTNb8+kg+Iw/gxTRjfi+WIM3lMTqmz18GUjDYFLkKa
GkIAZyxJIN1HDUP2h+RJwSWQ2sZbURfjAsNU+XwcjOAqMZqKWgB0B1ZLwrQobVC5eptBdwBndznn
Wvk+LrMLyFm6jQu9KWw3cZ+AN30DyoJLTYceJqiLINIiax11j7iiE/hToE+J/UfXL7a8AkhEYOQh
YgO/qK/rnda6kZvJ5mJHXNZdPbyVJuu6bZySg2TPKqX06geMcjURem3anuQUs6m+qMg53CoAbkPo
geUtPORGSYpywd+zdfyrPh+MhK/BOLFDvJO563h24TKefVNAKIgYCYQtmjCzMdxxPP3iAw1nihJH
fElsWjc+3/HpFxnsnFiU3XSYh0Kbrs61f+JwG6KJpBW5i+VO+I98sTrrqzSRSg1o4gLmlo4SioOk
uhgMCsELASW+xatcbJEfGbjOfs+gUjEjh/b4/LEQAPa6bmB64B92ahlJOSvXAMgUBv37pvpUAjJy
aqHu/OAVHJHnfsTdhGYzI/KzEmnzzZyH6HrA5nWhkXcmnIkcAu1PscObnOydCl9QeOZC8BfQyM+s
E0qY5dMB9eHGtdSK777L8Bi+v9bWitc5DJ2l7dkuV3vqNap2jMpI1xAEHhvNrsZJOS4ZUQK+Sm1k
YiDmUZnb4aMhxxQJ3i2lGLPhzkOKYX07AZepxCaafW1C5ByGmbG19Jheq3+QFyIKzt7KWdO14q+C
A442+N/CdDoo11fep/B625fvFZ0rXPWAEyV46szPlpYfsZe3wCiWJXkUZJiwV/PCUrxDdM92bJbt
dz2CArbwPf2UuW6GE0aAyz3pTHqoFCW0HnMLUujZ4NnsLIvNw33TPu1JryO2jdb4bv1gqQwPuqvW
t8tuYw4ZQ/QjSzUGuh1rH+qVvwCpvWc7CCRe18MqlUqB7c4YnwreSxLlMdmpD8moPC6SUDIIlc2B
hs1lf9C0gZbh1zGy1h7ojZu4PZl3EaZHi5SzBUWZgXXvX7wpAyHcFcNa/6hV0aciw3frqlf+pKyj
0rSkW4MKdqdXd6ovyqwhnb9YNs7tqAT5nxprtqupdKgU4+j0K7IFyW4K3+Rldf23AY6qHmkIZ8rg
lI+T/QshRmfigpx+633nLPm0MXL3JY5boZfnjuOPSA6Ca6P1x4cKJg9ILSEpYQWbDueoQcDpaRm2
3SNU4PIDk3dttL8mrDNiLFvlyz2PmDEHUkI6msDhDPUaTJuojxUXlDIFLL9NQ02m4RImGRmKrqB/
V5l5Y4h2dRb7CYr20SSnYOdqSqp3o7ZVWxZIuUsSceMchcM+ol/yaMOzjhGhkDxe9praRHahI63V
opwSPqBstzlro6PrT9xQPknEPIlqd6ir9k1fd9diiODhTo0ve+gnviSVKqWnwtVOkGxwyJrfyv3w
Scck4PvvkyL1iwKl8/ZGNslkwg+NuDD59DHuBRGNc39pS5/hwB+5od1eGtKSfVZuKVSfXMeRsqiW
dQxaNm8yzNZ0KgkpScg+1yMOqXQtpZ3lL9VhjM15aYFI+ZTJYd6NbekH710LtuV71UL5apQH0Rfw
CPiw2LnuYgZ2nYTdG+GaUdKkbancX/2CA8NCBjqLopZHVkIlCgty4LtWUMaRcmyK8owp2Ry9+BSc
B5WyAvpwA9UPyd/rGlUhh/8r0R+K0H2MQauZCCMdbHE6uC51HUBzHbJSRCu1EluvYeEvWSM5gDb2
F7f1ROlwbFs0CDcu5JGdcRBQh/5xypOsJTUxywm2J3/BklX91goErM7CkXVo9NGWO1DjXlMfN5NU
UFGEekVTDQo29Fgv4/Wc60amVTm0x4ztYAN0j+ueCMqesQR2vZCUin9uJ0elKE28enqdE6tU68V8
JxrdkPVYpwAlH89Ed2iK/NH+/JRVsWnQ01EaBvV9emFlaf7jAXmCDmjTyb8J/NNfGdHmVsTihlUn
3J5y7bXJP3rhkADYzjXPWjr3kbnyc8gpeMR46D4Y4KGoE+YtwM630M1D2R5VLDkdcrFd1GYo3ryN
dYvA1xfhFD//pSsI5NalukMPAi6emigi14nBEIS0w14tbcawPGnkZBTED2Q8M+C4u4N6+5OGGp8o
p3fPbSIbE253onYyy+zMMOCtHssslVvmkJn1el3XyTBmxN3Cp8ssM8yGPKwnipHZj21lDh1HyKzN
Zkp9hafFF7YIDIpRvBiSpL3ebhNFEF60qb1ZVWcaIbYno68yAY+/Usbegs3vfocYSTVbmApcs6K9
Lmj+K5I1gKfYJrZJk6l13WPVRP8P6hnex+vqnAxAB17vgXVT1btqu8RovqPKh49B2wLKH4w+4CeG
TlGfIvD9H2t5ZeinQCM/z8T/h2bG7o/uuwjGoNcWwdSekFgchJLBevcTzc2ubNJDmqsq2Ah2EN0X
MoYGMLklR9RQM2NWBcmyuHxpA35TcoKg5sVzYQkv2icecY5BvOL3mIyjfZuJKQv5Si0lv52MaRhI
ojIz0b839TrRVoVvj6C6w+7UXyvoQiQVsI1xrhZ3KUAHV1ca3g9HZRfEXzh1avpgHGUPNFmXq5yj
ajHblAmi7PpCd5ySBBjjpSPVr7flGasX0PqbfE8GqsHarVsv1IBE3VKwNxCBO0zqXqt9tfmO9f6V
oz7vWeSEqchCIOZR77ZgOuki1RqJFuwgwvOtAGPkY6ETuCB80L5OOy1K3lXeRPB+oQu271MVdymU
AIXuqmYqmL2J7FqSalHBe7n21l/CJnxQ+FzJIJiaPBjE8cO/5USHQ1/mI0Ot6iLlKoKwhnO+xB/q
KmluqhtSQ6ZXLzl2eiGLJK0xnGrD7HfFBTONOuKIyG+SgE2xpOWm1vz7pPYoGB53XH1wrIufI1o3
/WpOQxt5iLF/aEU8a049CBX/YxaFER/vsNuQ29KiN+16xUa8pCIJ6WwjDpFbeVa7k2ypowrBeZDW
QE19dM5lzae92dl8J+t4PvjwGT08IBkwtCdH9+PCt08rW+yGpTLhDiK7vDNyzGlYb396Mt7pLI4X
XLwXjR6SjjikKvvIeg/WTfGe1wRGywkFNCkF8x+0YQg5iigVJrT3rjdoVUc9Qj/NOwEw3q8s4MeO
U+yi8YrozdApEB5fpzAodfAUybrSOTWlr62gYl6lP9KLzxsVzDaZUhcoWF64HnFfPQQabS6Rt7tZ
9/YWA8fK2hiBsmxCcW1KuK3XqW9soTwECUX9ewFfDMDt30uaA4kqGH+KHaKsiGBQrx1SYHlvZxKc
Ron3SLGEwM8vmXI0qvJNehdrcUCoXy+9RldA0+ir418kGQ/2JLrk6xCbFF5L6oyiUXl4J8u0vT28
NUscJM/j0Pczp0S4mKTaONhTAeuymWV+OKhhsjZSg7VNGWddCiBgDqqu1zUGPlZ7X8Ntib6JDEkU
niPmRTOQgHipWNYPFfisRGOTii5/4E/YOoU9T2pmqXsCJ9G3nCBy2P2p107U8I0UdkZ9mQq/l4fz
2QwmmPCUVUOHuDNVsYqJFxCPyEYnxQ5cqrwcRfdipHGZxaQxEg9l95P3+5rTIkNMGIYz9+RF4b6a
u4ZcJHdlTA1mRv0nedrmpd3ccBpbf2AOGO6DhUGxh7rkWqdKs5q9IziLB8hEANQxYQtaoDaQvbnH
NLjxN7fqtePM1ykspnN840qYlKVYrIbNjnOGe0cHkUd1VAroO2vkoX0gruATkq1Ua7KrG0JLXbHa
yYgS5gwIG36KEE7ZKgppOl1Pt5FzOwlAii6ZS6vd2r/oOAF8qfa+p+Mcy1Nl7wMYlWh5ufhgz7Eb
IFJB2mIQh3pHPUHuoDdlTjxKvJjmMOiNDa4gSxfYJKW2k6zjYhBIzsrw6RYl1p3B0JUVVdHV/EVq
S4Ab/BZIF4uvqpvR1D86XS5U/5/yppK7s6NCYNoTS6v4kYwIJ8QPJk3EnCnFBihuJE82KwDOOfPT
qXe+ywKQa4X0IHV70flzXIgIo2UHQBv361aMCZK0p5+wOZo2UpAO5Ri3u3FN5kWhHX5Cymxn2rLX
sRfMW9p7SMGG2Njac1CEPuoeD9DUpP9ouoIwO1eALO0D34FdLXSC+LIexVVW9XAJc+yxfTKtwK37
wktIGgrdQnebCNcx9NeUJ6NL9d7FQQmmekb8gWDURh0FwEUc+P/y6/3zH0xk991i+3mugcBVgMMp
vaGNIf67XbsTqOuVYAkeYOvKhMxJm12xOcUMuCN6cHaoTW/cCf8PZbt3A3kXUE/n91JEN9Dm6R/1
V/AVPJv3ebU0xyeILzWvwQ7QwtH41JvJKe/gviJOeWNcqWwko8awgb+QN1xT2kq9Xyeh/Sw2XNCO
6crxuJ2Gthq+QxifpL+PzXVKssdwBWCPVdnBl6BMtKcmBOo6ArXCE/3AfXxxXdn+wQ2izlTVukKl
xUdq5YyDE9peh5v9LHWkZxYjEWnzFbRAM0Ok19uVPF5obGn95w0psg+cTO925PQxN/XRLvvdATfn
OLf1fFLnUZmp+IFLgWbXsDEarGZai8fFFTsO4mk+WrbqCDuRBjWZoFLdGLxQRtAGCcDOb5bL3+yX
aN88If8dsCuYIxOvpf4ROzI/oXi8InKDz6nnnU5Ju8qmFTN1RMYFhck0ixcZI873kBy1fr9LzUbo
ScmSnX1wBreDi9wjfMwsbEQbXNoFSuTo/wKNAxm2/7Ai5/Ri5JwQXkE1TyLUATIV6qV3b3/1Ok8o
qCEltl/4PfCuUjcPS45PYFITi68qnY6B0ZneaAvnCa164zNrW7jsUJTlZJ4v7b2/v5TZaG+rk2n9
zdkRkTbRrLndWyWq6KGXtbm0COXzmKtl4cmIGtrLm35ZVS5vipWne8TUZTZjta84o+IP6BZl9i+v
PURFjbRrz+p3LZm/ApHh77e2Fhgz8p1UHaYNUh/4+b4euZ5eqbO2/6ug48lxefn9b5mtY7eRaTmt
Ej61NV5KqXK5Ng9d7DVrqLvpeHHXfhd7q9ls4iKFIJHtC/kUyfpfPcKbDDEbf7H45aG/YU90pRfJ
VzucBKI0Znp7anltpqtOS4P0lOzalGp+kVB7BXBJquu1ARNYMt5Z7zEEjCzqp0RAKg37nCVBMDt6
KJal8TZtX7eJvPhIXhMvo5gzz3WFnBh/2+HY7bKu++ME8V7gjZal9x7jPa76czJXNf77PL3cy4gD
pkArgmawl60esJHazWjOhCaI76JW0/MRvl68x64SpnCScRRFf5J11jYdyCh5udJETATVEhk+4O3B
cfTlh5PBkMuJkBiDEEmm0XrsXaO5P9LtgZMtPzPMq8udRPnS3AOPqN2QJHjis/cYZ1l42s0+UrTL
GsWXFJPofVhs3T1v4zdexWsJkoE5vRHR0YUZq/4Uc8P+/rEW2JRdAw0D0J5S5WqSMMtya7g+UhTa
eMyb3WRdlj0T9pHgCSSuBoQSGuWyOsLFLIfZzSEgzW4WPzwIT3EaBqgYA8MbcyDP/SlsUyOTFNmo
LVc7q5UuUljYdxlv/qtdW7UBaX9sJHDEsCbRh4OA2NbS9K0q8WFBUBC7SjTmeE8Sg+wAzZbdtiUV
NeIOWjVWPPkEUyvyxIMUIw9q3t7mJX/t85/LYfh46iFzedVflfNBxjZ3e36NFHBLiMG2CaGPOJeR
PloCBSgXaYx6owHCOojoawXp4je7CKS3cOPuFmBeYrDLzoGsf5fo79Y/ofYijsto6mzahCcC2Pkr
of5+uGzJWitbdxmbIIDQ9VWm1ImTju///EPUUHhG6hrn300Lyk3YikvOPv4zTu0FsQnPjCtlI05s
VdnzSeC4mGmDgt2QDqo5EWBYAkAy/7K4JwJlknmDNNR/z7tVw1HLS867Z+eKhQLdHGq5Wb8Dbxs/
R0VmOAcM2A/scF9BtmtQDsfbUy2TLaBbS3XULqfJ2xRWfKpLCmcg64uf9xqAV+xCiTSv5rDzwUuf
N5mztWXk5c1U9DXNVerQ4N+LI52eQXLg52xpIAaivXj66Fi96OYE6GKrVVaB924qTtcDGczV/nM0
0AYcGaSG8IBHyGLfoPBd3kZ8yKjuBoUAHfcxopWTyBkEL1iFJldtEsycjlNAwDFMNKqsaMh3IZO3
4FXtDPgsBCfVLhzJ8jHAZbkK8QUY7WdCoJckH9gIvmU43Pxt2Ubht8WnE4/Ws5xQAQcIU4k0RU1o
mVdFXeODx4CYhKSox6G6lduXGMxucQETmMimPTj4m0710fY1KfhG9UItu4MlD2dHiaeaBvA0VA31
pJNnIwXHM/aKWpVajlNOg4EZDrSl4LbTI/KTlM/RsF3rMXON6KabT3CGq+S8BWUKVB9YLjGYRvye
1dJrNYCb8aVCu+byRlk0HXZ7s9aaz5uNSQK8HunpbtUw2+aO2idETBX01wRAL8OJNSQv6OLZ6E/V
ogcqssg3kbkskhESQqgKJza9lglG2Mij2Nn2pRavJNREzJYfFU7TVBkh1NTyqdI+IcRMIaE9n7fY
bHr0glmD8xIkyxF7LugBwpBRMUCpb0jH7gZNEHFXqDOUWe4Naw8FezdBvANEKOLIZGEuTXOZUBYy
WsJ8PiDUCXpWzn6mEDhpqv0kSQUPLY2SN7QS7dSdOmlEFL75offNHrLN4/k8szOzLrjb3zNM9L6j
O9rrZATnfj4FoyGwBhrvfCljzW4qsLQ3bzJO/JzvqrB5CuM+IBxEgAcRxlIaP72P6bIpc+qRvOFC
mQtEanMxHdOUH+mQLq0rDJukN4juXy1b3WxZ0xtjKJ+DvVKQPLtQBwpPvnTooBsifCXKzDB60DR0
CAIT7ovJe39xoSSKBWCvej2Hh/OoeG3v3tj6RzS4c/jPDhetF0ucBAaiENR1VPLbOXyGWOEw5VoM
1Pgvs8Xj/gFTSRklUWQCM9nb0fzHEOnHy4iYMGs+5B0B81BUv26Swmp98X4IZwfpE2FNHU/zMmzl
i/r6R20RfzrO4puUMJ72TG3BuOhZns3qZB8+kylRMuDn4eYrQdr+rAYxLobWqZNMxRqa18HGE5jL
HlbPnb4uVcVPj90ufiBdOI+LG7JbALlWtHYTI0pAEexil9XQZffoq7y2bCxmTwYMpjEA+dT45A11
F0GUn/7bGnPOTBP6n2otGqyiHMWCALG8xTCHX+UYOt6krC9ErlArX8s2yPjrhCHCwLspj3tCPvu4
oCSViROJ8Yr3eUFwZh+zvZ92/2Z4IxZaSznLf9hu/GfApOUu0oLt1PepOv9svBEwh2qUaNaExR53
+lA33rqIleCOlYqDfLQ7IpWVZsCDHUqvf61OIPhImBRTs6nabYHqdX8BdX+ghRY5xipaHgS/JVji
rURNDG4HL1FzzEec76NOIB8GYZT15yVOGZT3Xs4zijkHRzt8p3nrL6JQZDt1nq8HkD56MALqkj+L
eA5cUI4uxqdFZjEfceMTtJ05F+ilWas3RmaXgB+bmC1FAfIrmbo9X8o1dYmIsdOOg3ZUvBAbGAh2
YJmqZCjunUCPoe47vsOG1JQ0L5479qk9wHD9u3WSCZW2MWfbWFDmWYycUHSClOJpq7Cn0ygcnDFH
K8ylVG0o03pJZZlDAt5+WmLgcXmy7P/9/Jv2Wqi3STgIWPKuepiuz1Y4z7Ig/TvSYLaLWayt2pDx
I5UbP7RtVYrizcC5fgpQ7qXsiwHAOO/S/EJxyMfQmnrsbeEcbiUcD9OVlyTcgHVRCnziA3ZvIK8o
6TTeQdnw8+PUh/vj/r+gP0LrZPJKpeXjjboQOXIy04kGjnvU7xFl2cdBYOuhDIQkiPKgAd5bo9wj
P30iAJHrqWHLoVifLxzl70fJOZazO3zzoxEP7qjKG+83GaOv5Yza/ezSedLYg4auRAvF78vd6pDy
LjJpB081GxQfOfGpA6kcurGFMRTaEwRwQQ/erXNOpobGeQQClPb3abbyuFJqDMCZW7OfdC0QUUcB
Y37jOZ3CdeOaRFHc60Og5er6dyf7+PeGuv8QkqW6+GHWaE0HnYo5a3S9TOeQTtw6mwqKsd3f4LxS
oiLOWvIDYQIv3uTNf1InlRP6T4CddKEh8ZDRKHjYB2fv8tCGNgCVPtyV583fsGeMMelgPvdapAvp
N3FFa8BYaw6plmeJj+N4cp1aiLwWzp6SmjSwfObqrtwM9d4dHhFFy25bwMgjYGM5T7eGWSBJXaK7
+nlBqgYnEg20t9oawSR5FtErM0vnKh5zzSo3RZEfB0Fsr0ggnhDa9b3yvKIRiRUas973o0cT38lp
ZTKA4H+UMtu7nN/R8GUbqaLtVimvVNLeYrNJ4JpdNMHaD/lV/5CRxbqGfTQopSyj3R+8u4SvEI4q
2oB/G4YOYK/CqJyUXDV3Y7whDNlN5JCMWM/CDqGuSScLkkiZlkfdWZHbsmoSwJAf6iFlfg87VjQE
91oL3Bm1zLuTUss/oxlVHXW3ZidPmc1Gv8zhC8GxeTcy/VCrofnZk2j0vJt0FF6TWjHrOF1e8nnz
NVHmifFN4JzLg0f0/9Qjd6OVSc8xy7BCvDDbDAhExoDLiwtiimkC/NsAC0iFU1ESd8dtLOcCB+yQ
y/n0dM+drZ0sznkAb7LvijAYppL3SpwRwmoua8MpdpCq0gBbk0+CvSTNKlg332IBaiv7Oet1RjyV
1rSABeHWBYve6L4oQv789vrdpJfyK2FSKT7ci0m8nT/RDBbC9ijFhGNPSRJwzcLgo38VFxQGcFum
04IxIxslNyn2UnhXPkazp/vKQswU86EJ15DjjQZChFbtyyDKxeW2oR7dOnHuapxdtkRxOYT+h7bm
Nuw3vCaP/Xu4emfQVdx9Laj5/Uhkzx8b0v9B+6WBg5Jv+LGcX/qa9AWX01YKdkecCeXAegf4zzAQ
Bk7a56crmFeIIGUrq5lqAsY5hF+zq9J4bd+ghwYYmnYo4gYd9txo0kWRDqeeKvHYt0O1sabw3IAO
Am341NgfS36M9SdqwtuDFlUy3R3wpAEX/rgTJLY2aVY4C9Z39IqSAhIzr1zhqmsmoug+ChzyAdcy
VcIxtP2e6meohpelRfoon2sCZpb8GTJmspsFRhrehxXEjS3mhrrcxkUZrOBalR/oSaKHHZVD7zyK
3POdDJumufWOh9fWxaWnTClPuVYgw+nnuYlfoolBz+3lfsHDdwZ9pyw7uPkLD5prjRyRTO3QYd6e
0wIaoF8wETc0s4Rt6DoQP4BrdgHzSElnFEmaBdU/gDNmhUzZpqgGnUCtjMF1ZwipmUSSX0KTjerB
dca+1B6zsnOuK1aJjHEBtQuD/21daLvAI+etWMKe6cvSfqB3qvsfFf/C2JLK4jJtNQZbjM7Lg5jb
0TZSXfiM9nzbxR4jgQ7DZW57ATYRWtdCTi7Cdx5cnfCNcP2mGBx3Vc9inhU33jpAoXE6myCLzvxA
FjNF1O4RTa2ktsp0R0X1PVCAs+bfV4DDzBu3VAIiBajqUD7dyegQ+59X5knUoxbiWJ6KVQqAPvEO
lo3cCuVEbc7t1f8PQHP1Kdf6PcnIHInD3XzYXoOkHveKTm71okFVrKhMbMd7AvRCMr7QHh2Gwz39
D9J8Vr07px0+wiCVEz/akZ8pEmj3VY/RxH7gRx0jjBvNcK+XrlpS2ZRp0sRAHbAdRxIGdgdpRHCL
63lx2ukLQXmIJWly9fzupfzG6+blzpkLLkvXMDbilAxtJsQR1E+VK6Bmtn+cO/xMVJf1532f3b3M
EHwwl6QxW19yz2qfUGN/c8gBkvn2sDOgc2qvRYdBYy/fTv0x4c99Cjx/x+fTEWhdoI3BdJadeMQM
AyAlj+8EFLKB0B7HNUBk89fEQwYBkhbWnBUucUuYNx3e1G/XiJ4cbOqa2pmwnMis3LTwvUdWTcLH
CLhe/ahLDBL7iW6l5iXb3kuXQPalZm8+bSIuxdnAdR9QfUM6mdt77Py0f46WitcpDHi7fqWtUOqF
bnaPMW2fOEJTQ0DaiCCfevN/SLJ1GYvwQBvOpP82gZxc6KPgxd/fKjV7EJIFtrDHS9l2148hHDmg
/z6stCMEObRWbpxv2WeDYfvgM8rCYkJnU7VMG2BT9IituOORIyYOCEIuEqB33J5kgjzL+h8Lxjc+
L4bFgBv/DRBxGJnyp9DMHgMsmTGqK97FpsIwDnqjVwTd3x2bs0NCT4SAcczTFN7Y2vGXHmhO2we0
0xa+JJAbeKS8arT4v18OC4/qyYA7ev9Enc/sQ8qDUVk3yG/BF6c7LZGIDIfhBtY1mSnvtvtnfbyl
JIvkM4aJii9bav6tW2C7VPUYk3sib0nXDpAbTe0oqKvafWzp4S4c1MXs3s7iuY2+lsVxnQRysJy1
xGcCXN01eoZ+EzFzrig0t5bkhCClErZoF+DoZ5WHRVi2/PpPhafvKProKZePGc8VviNgYcWvk3RC
3QvjQGFg678idQQI8Bb/o6u/ZhYbYRWlFqi6ZZ+TllvjVCuMqgELwU2N4PGTbScCbeiQ/OMClRSA
pZuv/AyXmPGjPhhvj1U6Z5bUeodoogs7n+zN8IaJZ0xN798aEcXZfh9jEimA5Xm83s7226K/rcA5
gXn8+H8LR+0N2xjQWTnkptAdswN6hPka4uEb1oWxKl9L6ilLAB6WaM7QuJU1C0XWkes5vXEuGmZO
PTAIS9WLvblyIbfq6OdJFtEXiXgZCmZtwIzCYqwWQ4zBnGeb9dIvNevutJ5uFVrbduMQICOaMT+C
eMZHuAnkg2ViL7nt1JaEZmFJdSN59+tEJLl9QZElssdgrzlZH7eTSClA+UxSLNDGjB9chXgWaUFH
bI3uUepMKMLdZEb+XHA9mjduELp/dtwUQHcgZN5m+ALaSe1zm1MVMcwSUPkamT614XFs9NYs8egZ
5k4t+M8FJO9XvpuJ+rkrDxzF8COU3x9oFPBh3O8HP/443B21slbxGVU2rC+FFzVOpaRvSPKQ0nNr
ay7oHlpq3wBGZuSc9+A9yzzH5OXASLeH6fJKZJM4TStuXAOofPDrQwDL5FWyAbdWFW334H6C4Y8/
WEGVwJob53ohgrvczTV0wdVn9A3Yz3naUWnHqd372oWpITsBo4pRBC1u/Qi4/vDyLWQ8nH9Gg4QG
J5+TU6v7Dvo7zqzauuIbZfak2mW1PnZO8BjgTRjrimnPkEIExUAmwoMdKMGeCYOesYsf24kRn9J5
02M+FRSl4WzH2gdqZX1GcOTESbKdNRJ9BA+60N+nSHCcyXcv+a0t6EHP/i6V3Z98lXMJl0ue/HEV
NV1YHpy/H0W7BJSBGTT2xAGnpiiyCYQoBMzGSm/vLQsEvoNWs8UsvUCynUvsEsSCJfsAgavXsdDz
EOo9Za8glAvV5S++ozb5TxGUgvIVlOZI6ghUlceiwdNT44Cvz8iqvog/kqbLO8bNV5QIAGZuEQ8v
ua+pLWrjct6p3Zn/0xiEiQtJbZTg2+QEz1lVBukzqOwNqlNvrpr751msRmHZCjo3pNEsLV33Gi9d
Fa8XwezAn6DJ70YsnENc9/Ceh/YqZH3PVl/8aWSu11/fBuheXdqGiKrq4f1o/KhXX2Cw8EWZxnhw
SJAKZBEYeRZfkGSXKDGV4TmfWw6M0ZxihoMHZ50eTf8x2wFk1Sx1UrlsSaqNGNXI/vs+hSsFW3B0
BkJSW7e9XD6H5TQtstCH8iBUQx5bnnxMZgdHKVhqtiCmDJq13HyCEOQwbnaqNL06zUPcBDJu+/y+
b+Glxl/3G1txQODk/UXO6Jphk+RDgQe05HFecR5rjm5iYZn8lvTL6UIJzUW0BQkMk0k56VvdjPWR
zr96X6wtaiBuJcVW9undkyvngxue+YoQlqp58v9fiaZsUigr2ti0R4TuACXHjYq2GPpDJxI/oukX
5L1YCqlnlMjwSALmIFC6bB38Yy5wwwkcK3MGBG5l+ZUfus3vrWNJ2D9EdF/L1hg00BFlsdpYnnAR
bDn8BmddIe0vN6ngymQMYC4tVtujZzB7G7SWX7i3ZG/bdwmGgb2XD6RFpbtdXMExcSGBVoYh2PjI
SEB7XKr08dmPa6Xtc/Ye1vi3xM148hzTSj7vpg/q2PICzn8wgVXshQZwsNuffa/jvXjwPmDsEP4n
2LCh6t6idx9cWRgeO/XtTlxlSYdvb7TmYr3t0Ve1uEo+dhpX8exxRv52HD33D9rnsRfTkB6djFFk
93hYhmwQlvA8h2zckwcfoRf5eCuqzdNfSbtY/TAZgmnOfSJbZtLkm/4mg8H3ntHreZSoFe9hS9yk
6+chqwlH9go80sTbBIij8Esc8uKDuBbQwY//tBE0m02MqDHEXhxTsl2NCLVmYafOcAHaukBOTMrW
eYtKr89IdhY2lkIoIhXAspv6bV5uoEac6HbEqwfDABA1OBmdTYcA9CUpEnwRaImN3xqklwv0myCG
b/Pf196oTw2xZJF5L/JsRIFW9JHgWD29duooX57k0VhoFex6V/m7mNbhYfCyCQYqhCEt1cyW6JH4
YpoP8nFIC7NZMqfYNRpRMnuUWKia4rthaL9ENzKePMgNJ6AhCX/U3t9StDJV1E84ZhNbcAK3o4j1
8RUA1UEL27fGQWJ+PgXZiXSvFh3w2oGEoD9M39gmLbp4uIJQLIqcYDKj5D0VPOKlgIxYXRRbM+LB
5cZMqTgzs+tmLIiUuw2vS+Q2qtjy9E5cg7nYjHZV+7kuhZtJFqZWc/+LKZudrjB+MfJCiTiyO6yC
neSw+UT0Kdun5XAXImPXnTPXP0bdbaL/QxKiBMRe+FXSrNNOXzIu2/uMK7T47cZ+ikWRVNUotEgp
GloYylVd2dsOMI5DQtZZ2UjV4vxRgbpNSVRGdFCKlf3rU1onn3pUjtV7rmYLG2WdRgqSSj3i4d8c
De44vR7s0dYmkldryEY9gz4JObBFHBM1ZAe8ja1sHd12tZ5O6Nq/k1HRzZNErKzw1Euz3mZWdYAX
3d27dx3Jx+kKLPWhGhgto6vGxHaEKVLIW074/1M0aGa56TeQfLkZhJR2GTpeIYrpGT+HAEBy87eC
eYWrqpBG6i3JALTSC2HVSw9A4/CCmEMKXyivWt7nTf8gVVVp4nrdQYYK1DFTp/hfzGEtYyM9+lBp
hWe579jNcU/N8O4hPL04L27Gg1ririz+/t7JywYtZyLw1erw0PPbQYVteUiZEviphliQVhCewsg4
Cms0JW3PT7jhjuQOGta+boc7xfjlOaXRDzCQAEMyzird0Ja1TzwxpgGfLa2C2HBx9iN68Uww9mQN
LZJJ+n7YP2iXFbSqpLznMkoSHDfjWUZ9M/EpQn/Fo7vdvzxmbcQoet8FAGHgV18PAGW1LIsH5wVQ
tKCmsLZQjIoJitChW91k1AF+mH4qBUt8uRcLM5BsRlzfViJqxAMkzLsaLAC7mCGOrjyp4Z6RdFaq
DDwk18E2n6loh5xeMqPKgr4eRCyM6SHrTzsp4B9h7DTlUh6VPTrGF0sZkFRmXXVrCRgyaZi2vAoX
CfMZ8B/WxJglq9jRCuh1dSZXF/w/HrE6AFoG5C5+pZ9jcHb2TtH4EXGn9I84DFQjSYacWRAiehgJ
pjpLrOfZ15WOXgK5Hu0VBull86qMufREeKEkjI4J84Mz79vqfLuQXPoKkVx+Hb0EGOMOzJuKFxZ6
Y5RG9T69fU+J62/V/AojAkxwGb/4FgHCVVz5oEFcvepKIGOHlgq097da/ybxYKUQtlCj6ZNrjauO
KTJG/gR/+XqUQ5+RyIs4y3aqWUFVxBrvr21tE32KlbXifUbSvZkmk+J0rgM1xv+CnVylecexAXpF
1L8MLlrI9rQMP5jvBarCs9PZMlCAPjiNXJxcPUCBYx6r96q1WE7JwSrcDAxKXIBYUqXbKs99f5F0
leWnZfXVQ2GEmm7G0ydXMnWpC1p/Yez8PYVPqHNWPj7YRnJcGFPm46uz/ZgvdAGtWtDwZyZAK8kU
lBjKS4y7g8dFtJfIY/B0ycLcinSVJZUwK5VpMAM6OPk2FkOqEVQd3RC3H/OqMNUDiVlHNTgnA+SR
4VckiMgHgRhlECW1Wg7edT7Lbaykvrp1XrrDP1Z058G8ol01np1IZw4iHrgpUCYa6VDIChe9AKyX
+pNnJDs1GtppzKil6XE8oCsIG2xyFnKDFy1B6NN00EF8sXL7IqR7/YjgpUoG71b2XLqx9Rf7Oplg
IrxpYVA4treBlcBFnR41dENyg0+SzJkCl4WicXtp3kJkq613/1MSSKfVkjEVa+zH+QwbrPRvLOCg
FB1F1hNRn/vetb+QEoUvZJB2gY66oeA9XMSXp3bGNhlvcTOL7pqr0UFpZRWR/H+mPrIPDQ0SCDu+
/Qbn6+Co50flvWBXpqdT1FjY+NdskUEM+XGRbeOjwJdyFggC1k5pIafu9y/NTGrk+idhljmm/Wuo
D3TKUOBa4yxegfEbrLApy13yrPRSZNn7Duyi1b/l7qKGX0bpoIYLU0b+X7IdoKNYgphPxkxs1pRm
lRwJsxpYhZ60d/gZAWOJb4SkhaISqKfzzt/xui5AxYHC5UVLESWETPdG9MlDqtpwlcssJwhwOOIu
mJH1ixNEF+fZo+JrrcSxsXfdDEH82kzcv0psQFeHNN2L6Yw3HSMPzijiGpclNiJ7Z2TLe1rN6rhu
CSq9Ooezpv/3//mJUoj/h9vA4BzOBegOnPc3g3fvrbqPu/IyWYWyeSHXtjfzuj/nnL1tkczhoe3p
MB+nRnF1yaxwgRt/EaBnLPkz6MoiI3tEvKe2VyCGidolReuV/wVy45sJIb5R2pPu8cjqVGkjU18J
rP5DuPO0uqNHAYlfvooQhXZLqb+GZ9ePy8QhuNWZu4cmCn8XF9+AQcDHDVXUy5bOZBB7d9/+K+MW
FDmfO1RRcKDkZBItNuQkM8a8VYQ46tZiogJEN/+nFhRKe/JS9crlEerjaqTZnx6l0qvVggbiIa6n
O7e9aR03whYzxlq8OOvNBSbGYPiiWyR9OLXZLL4/c/qR9cRu90zGVCSnshunns1LXJpYVRvAlMe+
440H97RfzHUoYAdAHqCVSl6NYpbt71obVoi7eQlQMbDsVLskDTJKrb/TSX4ThVMecyhpHbndEcas
LwuNQxw3x+UE9cplKJOtycL0S051jUCU7RHkQmF8Fe1D9o2YynP4dd7fiHuQJNgRLEsHnjFTMpbG
MzBWHIlVU+5s3Shns+Q9ybDDcqVNybxBIJmk5/n16uX7GzRNdqRWlxjtGtTAyr7nocndGuWt7zCN
Codxx616bWinF5RCLm7x5GkduRmvHLi2gCUuLw/vqe7dq5hhcl5a2XWgolCFuj0nn4TuscaLvVXn
i+fiqPqVS87B9m0l4osYEX8w98c7VOaxB8pjdxeqR/G9qfOS8obVc0JY/AC9QXLEF1X+6TBYdrQm
h3TBTAgZEzC5MNdoplYMonWA8PBebaZUuELZsy8iEmtMXBBZZR5Ary+PLUm1zbTu9iDVLrK10Uff
tU/b3gTjtAL/dNrLnt+69Xk8NUlz1T1XEC/Pbyjpqh4ExXqCh57HXFYW4/F0RDlO72W49Nx5I0hn
j/3HYGHruoTHJAJAbwFA7c1y1eAnm1aK1nY4EDHogJFXqF+3SU4ER1pM5VwCKRXUpM5p55MOIfoE
nGNnL9eVmCMFnb45ndst2o4WKNhz1902c3DwXUx6elgfV+Gx+8wj5NA3QDj6UO9XVtEx4a/b+7ay
0r4A0Ra3Kw/EDyQMdwkbiUdEFgNCjXSs5O5dnsve50vmJoVxLS0o6azTFLAm/mRycqd/irsoZAVx
eF/XiDg20/sKZhZ0axfRVB0/mHQvyxr7jsDNEK1NJBdoNmPSydQX24xC2BdeH1axrMeba/Lw/av7
f9WsSSK1wYddqOtANLjaxv4kQV7ez1/ev/B5uQK0j+VwoN9VDpxHisK+NfG2M2hHuy1xOqUTdbwl
bsDJ1kjN3RV2z8U1Opse2AARBffITCOCNTo+sucTbSivyhBNXLX1DaPWR3qt2OJAs+p9NaloVoqc
nLUMHj78Cc9XyMpNT39yWQVNjzbUpGAlCES0VWZaDorwDnXfpqtbxwytL5lxJOzU8O+6H/qud5et
E+cGLLkv48dQ8BWaZG2enweTMpLaIiJGufqQu1/65a2jtCPKP1Mo/Vtgm0RlmeoSHfKGr5u9gije
V0OqlIib9k0KcjCiYzRQdcLPXrir63T9lrqH+n3VAA8kz/Rfvsu8F2EA+1hKehiQ4NS+b2Zjl+Nv
2H3tSLTFxtBYIx4TgfuPKhOtqdBZAAenvXjCE8acegEUgkPBAdaako0EIf9Yzgm/j1wpDplOujZK
EvNjRFntZLqlg2ksMvPiiNcIvmcXsONdHa2/LqR7kG7dkRIcunta3DR0qulQzrQVL3fePZtrjwmn
bhdw1kUAaoJHl8nW8sLFqO3AiAaeAwZtcpsJxA++82cB8A14N9arQalkvivd1J8ZNQfFxdIOTYIg
Hv3R9WIwUncCBHLUWN5ISsAd0Hrbne+VaU+uLIYymyrkWgHBWOzZObvXuz6C2xYWe3AR/Qq2p8gL
3xuC4jN+xGJvkFREGW8yV2j5jr6qxfns3zqN25Rbul5aYbM0Zz9Cl+OAkhGJLLVNIYABwnxEAq/O
KYJQ9mE5DKVqimb1IizqUJSRYk0fkszn/PHqV54EkwSwgVLv2cOkVudlq/YmG+2Y6ynxTxauA9/o
d/QDU6OsXIVWpsJnRhbKWLcPWbc5ix7Jtztq/6SjVzF7oK6iYYAM5M46AIQ9O/LsYuuYkkzCZ/R/
XGkn14IzQzOu8AQpMqpDtuEaT8mV6RQSNLafsry0kpdfNGGp0sl6FJWgc3BwKiMBoJBC3FYpXW32
FCVXj5jIXnO7tAEet1El/4EGEDTD6MkdouAm3coWQF8tJg0Z0hs7IzLkYALEaxJ0trM9Rdu1MJ7o
JXDL7y159LAyULaWQJU/njHyoMNwJi9uC2zKl/5HWi+TPgVkKCF66aXrIhYYPm+hgXAKHfWQJshy
JJUe5l2e+9IOSPN1AjFDu054U8xkz9r3dN6W2RK40aU/+Rwv3FrgzNd7nGwIiAsYcIodOsU03xCV
aFKa6sfExSBEFwzCA+5f1ve7S1PGonPGd6v97MAaMDJVgFtzscOAGyR+2qVI3R8g/H7Xmoyl4HbG
4RS7EzKzTS2FxMhGRXm+6RCndz8YBXsnpY26PYBSjq1gqd1K09WDte1Qrkz3gnOYXmG2ibrcX61Y
jYHNss4xx0NYgJQYgbrrAekD1J7OwpctQMNvD35bvrQHoEsa4JUfjHYKTZCo7rmhleKrqpviK0aH
iQJAfyp47VFj3IsBwvbgW6C+sX3TyJcm9XCLC36FoGlbDB5c+5upFM6dEDmAiT2zHfy3tFIEak7G
wU56xldHXQKPoV3N0HVqaVtEKcWtI61eyVEfr6wy/iMGgj6vSwLaJsyVnMLN36htXduDI/ZzL+5z
ma79fRKgofbpTMxBVWS5qKEIaFBVJPEPCfUXLffh00rDreNM8pd0t0vAZlcellzgOk8DMIK2EOAO
n6EoripInR8nA2ozcgnLPXTZd0xTNO+ovbcsDbzdb3Jv+9kikP1hvQ5mLPoXcGbIAUbn921MI3Ao
z504v7MCswrfk+yfqcND+HZFM/3ctJuqrBru/9TgCExfjVXaC4wu5h0KPGZZUZJVV821yEnuLHEZ
mcznUA7PK/++A9KByUY3YfvouMPgDDLryagaQnnUz5FflrQrISgmSkiujEJFCsesbU8g1dhlTXCb
m+3sokD51I2gS3bxY2ezx2f+1B4Q8Jqj9dIsgDiMiIYfH6sKUaFBH3K1M5oG3tfWhxCxAN5h0R7g
lSbgyVCouz56nS21xa45YFHR4mKGs48dFqT4ZyJJyU5+lKLjH8D26yVFo4FFLEHb5Ct3ffgcybWA
bI8Hj7g9z5iFmp4SShAlLgv5NjySPEgt8/22D1v+XIi2MYOmwHqLYHPC1dj/CUGmp6ajz+Vax4Q9
ytAk085H8WPUMfQ5G/grhxQAMy/9nCdQI7X4hruessjLc3wj2TR2eciz16wfxtM/cD8ANFboKCDv
ugvpH4Bdqvg7JkmzVycptzzOame+Hre+XxF+xS7TKvLj4cYGkcrhD0xNr4S3ArXn0i/A2Rv6I7mU
DhvVFnpXo+y1Fm2SLx7okRm8EZL0nha8UcPN/fkXtMdkHRU110lMDG/Nla6YRZBze/zxoHJHFZQc
99WkMeMBgEYPzSYYCr6SQq96mkjA66axPEnr0VL1lrGaEHdN4Y5XPrimZytPFZMOPj6UIiAglx8f
wOYxhykT9GhZ/lfS7IZhB6IEuxFpiGUODrg/DuZk6a/eZTBpe5yKq0AfDhEsfzM7GoPwWxBhUXtt
iBrFnG56f3PpVnMLrRD0YOoN7tauCfs4D2ntjp7tpvdUt1RWhuxPgb7uot2ZD7efvnPAYdzqy/J2
ERb6Lz51kK3J2uEboHgezwh+HSqVcMXpzyXIY2r7RwVlGZFvYyx8J+HhnhsDEnR8J82jjs6L61WN
ySqBX5AldnWD02E/d82/pldo7sxBQ06ZBIx6v/ggI3eGOsX7wteoLt5TOu36y7zQXS8oHd7fpA8o
2X0fuEsh9z0nv0GF2YTm6I5NHmSMNmRxRPVnsTiYje1mWMYic4Drw5nI3yth/qEYjw4hm/T5Vksc
H5/O0ZS7T/6EuWgiP8bD4dHyEurisn3FpULYWxsil2nIaYQR5ZCdL0aM7DD1kMPOGD+tXinhhU/u
n2MEZI2RnTIp5A2Lk4xL29i6p4t0r6gcKm5PEhuRrZ8QYdMmTdrz5XwAURiN97gFrF14YXlItVp7
Sy5/gCp4gnWMup68fTyzRnfy/LfriuIFEvZzrzJ1MabGpq8jYqWQ4MpppAADgY9CLvFBE8AxLv0g
8YUBFwi1p3FnFGEED2jOVhP7QvEZ40lvDwzEWj/u81nRJLvptaZ9DmVMSqoZaqrNQO7cPO7JljlR
daNdMaNF0P0aAjCt/ozoXFmrwkX2PdYGh1acAW0dJ+5ikLSfQQn7Si8JmTks1IwYmFFwcIwRzOq5
zju2vPGrBBPys2s/XKVqjmPz3DRsQT0YNzJLJBfTW9BVRgDPiw4JtPZ4hniS3qYvn1JwzNmJjXGv
B878+Ex38IT/MyabI9LmfjOTwmrg0xiU0ajxu+yjuUItV97+vSz25G40awUZ9daUiLthl8XeFyuk
jHLotbBOgblX00Y7T4XwnYz9IOBJtbPFgRqr5oeTMrrIvsKvOgCIBfpEPgg8iCnHJ/+SdWDgjvqc
tmbsAbz8WM5qcLyhryMsPJi70POoqewBe8wa/RH8bPj2VhKAjr82PCVd8CaM30gHLkaF55nJ8CyH
2NrZDAdr59gNSRpNgm+MNOwnf7Oijd1wjK7mZgKo8cnMIz78qYi2HcH9QDVDYH3N5Oz7xPpU/ZWV
U4ZZVYLkBxd4Z1FeMy2IJPwC7EDQvR6sH/b3G85bLrkbOpbq615s+3Ba7MHKF/VSeiVqR1T9S0ey
3e8356zwTAMnRz53BjOEA2wJB3CKX/qekQAFo3VMlNzvDK/rkzCE9T89aDqkreQAz2vlSU1mRna1
qrCf32MfsvRyNXD0bEUZeDxUAO1NG/QZq6t4b3uIwNh1HI+mMgmvVyi2dK0uf4aU8bwKSxEH6Vva
bgstB0UhVNd3+RjEnPC0T3asgj8t8nrDuDjHuv03Vg7ohWRAvGziNZyUndFFq0PUI3Kadjwi+D99
xbBjmu0oyzTsl8fSTmQYihwA1wWOI/5xdFcvOJUoa3TOQEiPYwMzvxdBJz2Q4UelyauFr+d+eMrE
KK4fYRAqIL48r9XK/pM80J8j24j8EXCpze6bT7577DdwGwn4a2/xiA15CWcfyDMyme3X9IhnNrj+
ZQ9xFE3ukklLp8g576SapxJgDeSQcYMw6SgMXqaJpThKdIVynKzK0+wFdoDKZUVz30C+9elpxBTS
fDR+N6wd/oBVeeUSGJzwWtdse61D2RY6aTadcTi1CRItKq8z+Mr+bnzNquOPhTsBeowBxrGIJEZA
2Ef0PgOAbZfnTPhNHGkkUerFVD2RUud3e7jqQafUjDnQH8215ILbX5ji1QELjwQOXoGIZYyjugxt
bRlR/2EHyyWUGoPIRJ5l8bLvORms1xU1AqlkyH3leGPd3PJ5TfXvLTckfAJFsqiyEQikf9wpgg0D
ZkmR0plQuNyxmh7OP5SzmbjWPA8NoC1RzK4U1NuE6fbPJMfO2KBvcesOiDllufq2X46LfVZ5AWiv
BKeGfwsM34bHbw4UmQfQM7WidfwezMEx7hlYhteesLJSu2PQLaNZfT0PTUZ3TLXzz0ZYyjC+XVKL
4QsTcEjorupTR2EHA+waopX39FllVf1tHRRSvp61T0e3q5EQfTNXPEb/GgI1dReSfGqRixg0261x
qHFuHgDankvEZj4XWP7yq4nM6VFmtWohglM+F3yl58kXB92TQndmVSDZh9WryV1R8VC1dFxnJCQL
yjC28PMSzrKVa7+2OppbMM8om3cvLTSb2MUZjyqdyAOfvNsT0a8/0az5zN6OK+zhYUk5D2Vs8meH
cYNCA2Os1DVBYhy/WDqzdRFPlCjhd2OW2WCx6nOFIeer/RkQib/ZyFIdYQEBnxZZ54lq2LVVFZQ2
qIjDO5FairiQGz20w8iniz2+y65TdbmGHFpuNBRmu/dg8vHdMJKn+zkOSVVGo4GxNm631uB2a07Y
AHaxzojNfhcmNL4SoSmbm2YfzrqxWD4cgzmhnZIpEi3D8TBGkhx598oM3Ih/1w1xYS0+wVFvuzDI
k9Ejtx9G5RQzbzuCfdOYBAdjcv/jl5tHWY6BkLvEjmQCi5xxEXo4GFFPPvormRHpK92kdCAUxZfN
z8NiFv8xg0k7miOQO6c1YOBqqzorF5t9o36ObQ9zmy8Q6hMXW53WlahuFTZSgBI6EJTP6oPmEOs/
qiJ63mYD3Y5OkZ13WnuzNpZYjQDvBa2TvsvKqUks4Mkfx+nUkiyApaccPfd2q3F7pVjsbAxErx0V
OOYygb4sbLMqHumOpIDeOB1931Oxjc/ZoafZrECKnq/PvjL9jZVUIah0KBUrsnnhUKGbbp0Smb1I
60x7gPzHpgN3FvH8DnkwEBkXn/XNqiXmiHnd9TIKv7gtdMWXUrtycrHCPkYaYV+2Og13LD8syjQa
15bL5/OZmeBiOiC5RNqN/aFgB9usSsEthfu/sk3ahnvHUM+bXHvdBTd+Vpcrvh5ZzWtRijJs2MLv
XH7YTwN2UNvYo9+rfQgPI/y56o6Mn2ejAXo1H2qAqde3anEZm2L1Z4GFKblq7pID9FOwF/hcxPx4
Fe7ssq2aZ9M33le32O5HcX3It+RkWZczFJSLYheZP5fedNNmKDXt0l70paGUAQKdjQvqt3I1+NW5
Dq/2gZswnDQdwtnYE072lSmetC+WfhY7629q8v/cDE60x8Lb0QkN5XqvvJf8Kj4dlB6zoI1IRP7c
SxGnnOV3YKU+yxEyVz3UaScUcR5eUHWmtZ9vwul2Cjue0M8/Nu9ft2CnQNFWZaM9UDmaymkfc36t
wFKALkqA+tZQKKCQTe/1tBnNe7GuK33Wqxs15QZ7YLKT3tcWhqTn9n7bvohavHK+GYBLS4ccBptK
1rHM4+3fy2J2Q2w1d1Mn+e8lWJx4G5R/lmLIL7FnpvHaV3au9Vp5SIT/N2Djzvx7cMJmUSQrV7mq
dPiXg1VkVfG2zyDcl9HctGgLOaQy8fvDRt5qNTs9T3TszegfpHB1YWA0c7NVwlL9jhbBMgzuNVp1
RURaG3J/Ot31+rUhHJGVUa2hjC3lPkEw4jzGWnScZ56ccBcws/nO96s+QTapJCLS6VSQ2SMT5vUY
NviL2T4h9FlqbHojcXJueN+KUNVqPASzc6L0vMIo570VDligUm75IMXTEAPXOv8T48q33G8CTbQl
z7+ane6rRVKQ1tgwwwrTaut+7RAliJPRy68/Xvh3WcF+qUu2m7Y8e7Ax38bekcyRDX7HlimTuAYz
wXALRnBexA1fb1AS/GmgcNqRWX63FAZrEem6lx0AImeI7gqYuNl/dH5ty6bQE27+o0v9F6OT46dd
is3oohBbMedtpcZLXTkbATr0x/dN7l5AE7/gZJd+9zzwT7gt0wRgb2AkmgqzuISN4mt33u/VElWJ
ItnOr1dH3pT71O0TOQCLQwBzvHz7PVgg2scQi3P+9thg/4Mpsa4cCnLiDbqkYVbJwVaRyicse1Ab
FTb7o2CtSEHzxOtu5ADKbk19rFkWdKd5sRFvVYQUxeT+mQiYIxibZriSi5dsSaZs8b9EdzoCr2Ay
nfkU4ddh2g/D6MMY2Cppf44BDrQWa2vXKCrXS57+D73tj3dGSzwKQFiKuzPABP7q9hfNgrB7JQy6
QLC5HOPD1Ula1kN7Qm89Ik2cPLR8ZPi0/yZXJj5/u0ntvWCSgdJpWPzp3x7PHszhcnqTFjayK21T
kiB7cnBfT5pT3V4kWy29aac7qJLVLiBzWOmNjT1+it10OPfpB9wM1mNZb2Ufc+m8j0Gd9jcfgfGP
siHW0PR/JF7pHCSOSQMmTqPNKWLSdwTlJaHsQVGUHAH/OcMO0i7nVyQ2RcACeEMRljdEQmIN6iwf
B/DAKPLxFBfVHnXKfWmbWiW6X/C0drDAwmUD/DB6pE5x+pBCNPyeRxcyN6fgTqNCR6A6vQwzolDH
W2DQKIK3aaOs6in3e9c6OtI27dqichSWsffyckTBlj37qW46XTsmDumOKR3y86cgsplFuH16YjVK
krKoaCcj7+BN+mv5fiYNPOdIDAsQ0t/1Vfjg3CQkRFPfqUvDSgawqy/HMp8ldTPFXutX6MWDuyJy
ymIouDCT53p3KgAyj+dII7VWdY90Av25X7loYNipDsWZCRZlSIjB880Uw5sYOcRnDGy7XD0suAwg
D3h3rxpruDa+6aKI53Ry9lFw11lPRJWBlOMlTzaQEO0urrwlb480yjd/3VnYO5P5bGjjk+9cgU/C
EAo4yzeP48ZK1mHmt1lLDR95b2FIYeNltull+fmXJIAFaQLgEOZsJC3NtxH48yjv7BYal0/8SjMj
rfs0vmad292uqpuNIyM675cVU0rGS7Vw0ATsKJlosrG+94Cr0QuIdLeqKgRaB3BrWxnUtcABjSGn
+rOs3geUiNv1uEYEiFUVVgZejn8DPzX14PgByXl+H7t8rDDFrPhvcvr2mgVpv6/XRtmIC6Cv8u5e
cTpkMiX1m5kXkSYZYANovk3Y9jnmTI4OQgWeVyUzpUBVK1GPLqpftZBBL0yRWjOrAjut2b9H75/s
6JdGhRnxMpJ48Kn1Lc70TqBysb26w6I1kJ7Y9F3B4Ja2xzoRXp9TOnPZL9sRXGiiRcaoR/mO5UNd
doZBv+mgjKhbi5YiVC6kKaPdFpY1zGprJC2nfvDdzHKylojU9vxMgL0ERXcLdwB7asuh2OSzxIHa
Btm0HOUJnMu5NBo45jq8zQoQht67tCg4UTFSMhThFno0f53t2SWXNV2tqap8fKIAT0HpsQlAr/ON
kmkYumK9mYvvY1vkTfhuJySiICBMlyxxjW46kdPq6HQ+Vkf9TeWLwg1vGN6S+6j+4zMcvSZXOtAU
phswQhblakOIDGQNaQZ+TZE2heoyItwV3G1YG3CM/39ZP/8PuLDODOr07M8zYbndmcY2rsCk8lUJ
sNO/ltBZ9dMGA7/gp7AJ14r8e5/zBNNt/j9SeDSRZpLSwUFNvlfi8pEQXZ2Lh4B0ViP9olFPqVaM
lzwjPlPq1wZQFIAtJc6L6+tOMTjFyvhb7g5//TrbuPFQ1DUi+JTKDwynEWrvf7bz9G+TWgZiM6yP
aL6bbG0B2FBAQHTMjpkS7lc3vDcKA7qj4sRe6wCpn0+f51wZNH1Lw1uXLD2n5OFAk6/AGixH5Bwv
tDEbLZ/6z0hVn9tjR6ZJDuzK9nh1I5M5CvYQUm7xjEJ5DQap3CTmhNLHLMsGKfMj4w/FFFL8U1eX
mSLb00K31rsrm/KTpMCNGYwxMZdFXnehkVSeHvzI7Vnaf2W1djRCTyosWcNBnxIxd2KdkZVc57iK
vyLitB4Xs3K+oPdQ8fiO5W6933VUWRNyz0iv+pMYmSKR20G4YW1lE6zE2pWbymO2QQuYutDkFObo
1Nk952qtRRPXSF1hYpJegpafF0dd1BVrmdyRHfNetGWw2E1rAPq94I9tKhrjaaaHeAOJZsdw41sp
yfUVuQ3ylVsT4vGUbNj9oDRievXoHEbAwn+BpFgeOl5BVTp4GtS9Q3zPAd6gtADedmaUD/mzuCEa
yfa4emwmJA72q4Vj3l52DfSnb4xyLgVMhWhnm90UJ5GtQIC4bfoOqwkE6RyV6caWwc+8BWVOe0cb
8vXDmWHQYn6RoaCK8cWDyEOwQfthrCEv7mvrZKQGDHR4J5YkkGSD8aqaWwZ6vTrbaeSb+yek0GHE
O9lpPUBeNakisT08jeozpcJFSIEfcuittzOGw1zEeFI9K3tLPuwJh4NxpZP3EFjnLQs4t2p5lzQ+
TiLrHeOH622ia8dJdXQHQwbhTOHhheQCLYYb2uCGVER7Cl8/grDX5XAgmDMl5sgIUt1ZhB/vfcUd
qwafI6MKnuQN1u6Oa2pNksz/wa/lAhONh4S49nSWt3EDJVUfIGLckFf99jVX5gxVh8oEljhjv+uP
QtZC0z/zFIBBJmHjCBjOfCwjzWAEYA0Glzuvyo5Fsz7SN3Ue+Gwbz2bzMw/So+sfFpSJJ4RZpFZE
rJIPn3544n9+hTSRjSB5cZnHIgtZnXNQ4Yzx6/HnD2taFBZFlJwBdx4KAL28Bm2foL1ekDXM7xGw
iq+d6FQRPi3eEY1r8Igytf/44E/PAAo6w+zzGJl+z4uHcSK5Vvy9jkRATtPIoK4xUaCWZg3fwRBy
hW23m5PDKtwv1syrKCp97nCotS5Q+45htce9dbxUm6t/rWOSBgmKrzV1MnmbmtycQq/T39WU5P7B
tX7cYdV3VWo6QTdTPDeq5bVmZp9LqM7T9F5QuERw/7ixg10ca7ySz8GZhrqO30vhrK7QSq7Ii9kC
kPKW15QwEC32Jair4cijRLX7y/vZjndetnEq2x5jObEeRpBjFObVYKkRMA8MHDazN7/QxsnJ7l1A
tBLUVrwZbKbfxEAIExxUDaSbEO0rBgm7BgFzovYGip1DKghV5BJjsWbalJpISBjg+gNN+cm88mv3
V0VO46R+zmNfviM546pdbfbB+5upsIUY6Ki/f33tGnxqz7TegpHOmDYNBs/WuuFcmbBiMpMa1kgQ
Khf8tW/D2J594M0QAeLsG/U/famCJ0AmQnVYQewSu4o6OhUI0wTrMo4fKSFUqwWgOLVmp9QqdGGj
0PMbnc6aEmIP7RKr5ARMvS0f57pDHBadjtbxHumO6fMz13fv3PZGyp4g7AlOKbyKNesqdsCxhS3f
BSjEbgf9BJcnVNgCone4Me0JeOWdYD7Ikdsh7DKC+LzdA6ygXEWT2AAVNN8tzYlnuoOdT3n3yJy1
8LjWlQoGE5Lt8xRZljoN4mvywLaez/C4e22tszta580dsKLpZ+Jrc8u9fxasoUH5MvatdOVpUMdZ
Mtudb9vVfs9V1dPgy3RsO93i0vpV7aC8T3dvBWQw1/tMRQmJmsyL+qfj4RXa/ngUzXVODBOEG74F
b2znzkqYKDqJwBoa1r471QEq9heR8m8eIV9AB81oolBQ4GlMLpkyf22E0Huv1AoeGD0b0OkZzTwe
rEhOVZedPWkJkpQLKaUo6Z/wEiffDh+LZU624M/wB4ew/kor5DkCBeDhDZYog31KdJsoTVz7Dba3
+hjfe3Foo56YiRdXYJyThncus1y4ECST2is69B1HV7AiGBqLWp79VRkrQsXCK7Q53dECU0yv3ax4
B7iMzbJ4AikGj8OrsrVdNj/WfH3kMZhr9IbptjCV04pBKuP7QpOwamFY1q/4G/E/SYBzU3YeRHlV
uIkzByirGojgkTUUDyIfecOAQPxVmwOj4wXV0Nt9y+aDA5B6dfeCKXvfFuI+nnJb9IIRvEVdzW9S
f1hVFgocV0NYShvwmwVlLgvemh59VGpjQe5KvicfQOxTToohThN/N16PqCDkWag1JkDPq9AgRxVH
IGVBSCUjp4aZoJyNOwq1cr7EGOsm4vmVxzyEfLsST11/B2aDqt1YRUKUgzxhPNQPY4PpnyUBLXSm
f8vQ1sDE7lR/HlZphyPJ1LXvDBGbZrDVakJ13EFZkCl8G9tCO3JWb8DQYBV+VfXJ4Cx5fA2+kbM1
bgMgISJVbQatlNlzBafywPSiHy8iW5b/ybrQjTlKsTNVaOxoTqjxQBkx0UofQp5xf64j6LIkvTCh
i/ZOTcxMyu6B+g11oHCWmJCuaqsfxacBvgGoz/u4q8bqer7yB5oJayz/uWFLKWx6HUcwwIlgSjEr
tS9LCs/uwN5UM0wj+93z+gYYhly1wxXYgjBvk5gO77Ca6pmy+JSl4KkXFmZgAnXoOouAk4Khl1GM
WaS99qKZiyLs7xQtUJebd/qkFuxo45DxKDSQ5/xZqqOFd+UZzq8wUuOHM9k8GWT0m63KQZknSHdY
Zop4CFKfFELHiT0U+c9ZXOdmzUp2FAYzD40jzB64SVQnsnKMc/uezj1mYDrCEIWNwvFTFyKR4bHU
LG5b7Q3z/XnYwVOesrNQs43fw3a4cExnp0AidVFCnK9IrWz9V/hlE7+oSaNXyGtc7o+bWD4dTr/w
sZQMps9C7rC/qE1TMOViWpexZ7IpkI+yeA4/h11SdrBmXMgimJQe9H6LflMbxFEZjgwam9zM49+2
nsyMh4r8e+0EQ43QfhgzRlB+LJbvZZzLeAw8R8KbqPN7tzM982w7O2M7a8/QkE0l9aameZOFmXfZ
5MJ47rWuhoM/zhiTPLSf3Tcuwq2WMiUJs9kIQiI7c9RttfF2wNnlMIAx2wy2mXx0rogEwT5SHzUn
VEHuCk3ZEq2MzOmahvgwa3vne8WgPJWdAbdifd+7yUVbHG/b4AE1lNP1RD/T0qHBghpgFyrf4bbM
wpfeSP7NVBLUVOArvldwUvaQLf9UcMXNKmEJOQHfNLlq1lPxI579VG61jVQfXJ34PIVVQ4iVmg1e
J474WzeysDRj0WosZxUX+uI+1FlwdfXbo/7dn8tWO99MY7OHQ14F5mt2kGj8C8074m6epwlDXHy3
UE2GqLSH8Tgg+2BIQ3z08okKhqtv4CaR1N7m/HWbbHbyz/Dbmv4qm5y1VADyLSug42qM+EVj1qHH
r/XLVMNFdj94RKaUrlNCjE4jYVP+a+GFwkr3B3sQmjNrSmY7TIpIgH+1hqmf92sXCKc3mppPSVo4
akY/Q7jCOdxqHC5SR79R6YsuAGHSPKPtwMUw5lRDMw/oYFmGBZS8KHYT0NaVcrA5+tJ8EvjPlH53
gQaXQnekazDZjOvBxaBks80C1P2I9wnrNTIGK50VgOm5qgxCUPn/m5yA7nX+P/ZbGscE0cg3qfJ5
CMl4abhBeaUzcWDvjeSKsBs8uNUWVU53PpvH4nKZesCJlNFvrV8OEmf1ms9JZYbrynPKhgueJlgI
YJ/W5trLQohgLWEdBoKkKxRjQ9jl51yvq8LLJMRzCpzSKoBOm/HV941+juE8/4WJ76NG9qu+Djir
apDQ5YdWLP+0hVlgyIyitdz1qbtoX7wB2LIRLng3IqCGoWXMupD5/r8NzfCcB4vZy/rhAkBDowjp
hiqyahzO8QZXQVtlv+Uc4xwm5pCkxgEOTzRTZfDeFh3BmUr803XkXShFGWi+1BdtpBP9MWv1Os3v
xNftezAYfsxu6LGr7krWgp8YKb4GycQZoqZyZRych9v7uT4aoVdfpMi0SSCCMsFfimMT1MVWr6wv
VwvxwCiqXqn2DfW9VEHVM+QFwNxaQMsGAVaq3+0fS+McSNKlhSBZeKTtmGD0jWnwmpyxtiG6S+Rs
nPm8v+t9BHSVxM49KLg2EUC3gAFzzN2SNUjrWIOUQ6Tzfhg5Jqx6xXtc7ebY6fHNsmvsNvLTGCax
FJxcBrtmc66y6tZM/Uzx6wRfdeMgDHMO1UsBeNhPc9y1zUQlBMAR7Hj3qH9XJhyf+oA963fAk7Hf
ZHRkCxpYdimbfOPIP2aoV4+uIAm9aYyUO+gEMYryZI7JvluwfVZiMJlH2oqt9Sr1J3Go3S16SAjH
Rt1m6fWQYedvTXjWJWv8/Aj3vxDBiKKPbkW3JHwKWowaHfRNuzLGIOwMdWX8gS/dlmcYzlWZTLny
V/j8ohHIz7xsdZZuLkZ4NQBT9ELE8Sw9eFnszgi3kItZZLNf4mIkGqZ6YOd8nb4yNyMJVkJ5eExu
GSCuL6oQy1jENbzdQM7ubYhtCFiugd53kfSMqNmGWrUaeXcmMbS4Dsp2WHE6rf/ejQBjndDcweYm
7IKdv5pNuvvrRXZvkOl8HKaasUOz7hkVjANDteMcjpS0J06u40PzuVvzR4A/JqWTgo+qkzxkSrUC
PxgJd6IiQ4mk4acgVPB+hYPvW4gpD2BoEusyGcT4Crz5TTKNJvhR8ycz+2jJlWwLoKeTZFCDcaQs
xLsY/WjRmN1mNKYH/bu0fBBc6eOV5gMdiRDZf+xpnhoKx3fP0MZBdaJWdbWGxbFICb7CGDTtw4cL
RWzcGLBfHuwNSOPoXaZPU0RqhFd3plPpiqVN9/nybFxPMxy3H5a7SjUoiLmqZ8lJiReGZZE6sZqT
I2/OCR151kzM4gZ+cRiEETCK5oXNenEcz17Fh6/KmebB8dCkuTLtJrMJsxx38FGh+Q7Qc4znHU7m
u93id/NdQukKpfgUx4A9WwSjOdZxVC5bZHRjUzpZH49jUxDwjMJgYDnbciQU7RP8VmWL3hSwZfi6
d/1Q4yYZx6VsxHSJSsKm6NUEnRgZBMwUol79O7ht+eNS74vqd1JT4jYjAlQfZedYTNHHdE2umFad
4GpTWWVSnOEhHA2TNFYzU2siTj/ckWh7wXC9BL3a1J/Pwt3zQmOcCDBNfVHg6WWiLSrcG3UKeM/P
4707K2vXctLk2EQYt1P0ZralaCx/5VfbGAGwwaLGOYIxvx1QRQTIZBQKpp1MnPgu2dFdFS/d3Ch6
nziyo2ILQYWprXOGpdH5++sPmWG2W70NS5Kqh9dAcPp9mswORI0gfyhinLEvVMp5eQXEqE3nRTRO
lvKyrJRhTJYVbY23hq5i/2uDlGZPvJvW/YX5pHVb+3Pb39dnIYV8CeL1oLAo4qwhYQznHPo0C8tY
y4lM0kJ6Jx0WpVYvjy+5L2JTnGOUkMFqX/knkYed8eRp2DiSgRIYC6oyWWnZlxRHFraGNDWAjOUA
YfDkzDKWvULSDfvDZklEdCXYySaTDS3XlDqJ30G83LVrLdD6gPDfbWZefz31iKU/GQBfOUlktu6l
o0buyQ392LTYl+GFJGBjEqoYNDuTH3iMh27MTJHwyKRiqcR4bQdHillgDMpPFJJnGDo7puDCfCgB
NZLR9QhOvuc/CB9+d4KgsU379tBm3rU1taUMx2dnpxiFx9cYbdAHnlPuYvFrFRs720pecJSR0u3q
MWq2ycijAmVCT1A5Rdfg6jcPT302gXIAhugQ4EHb5tUYQxT/ToEBjTih7OUFZqlNqzuBqnbjFaU6
o/M37jVftqjoKt3BaO/s4yVKCTcWPUlOI5yqc4oqV8DtT7447Vd+J94qwt08nrxUZKL9BhjLcoqK
PX2Y6f438PSn3L1vbvi8Vh4dapO083v1n2dObm0Ccnx//z8+I3S5yyrGdq45cb4FdpQ2mN1H7sb4
VhqAzw3yZePRfHRKwhlvwmeUSFnN4mHMjHvy65yWFnwNHMdwB91pN8rdbdOWXjN8sR/W/dxUDApO
GkbBAiDJc5CvAX97LIh69A7OHXyhium+3tHcu7VX85+i5UVaU2NXiXPJ80HXzsILTyJQXYaICIgk
R5GKJNMIELacaf7jC0bP1Hmr3tC9GGM3V3w6oQdDbvQlF0uKDX9bMrZaDgs8jjJIkOXLDEXAJzie
8gLklSB6LzhVCTROeA1SdSplIDCTOdWhFezOokyAWcJZoeKNgyR4B1uMWKefS81lHdUtXdxv1Asm
0XfC16WU8ngbotiOAdMYDCF7t4Z1CPgoJ9ywAurcgxygEtK4nJA5Gub/MLVI9dfFypfY3DKNUsPC
JsVssf2xt2NGAaBUYH8Jbe3yDD6mUhhqWNy/Gfg9zKM9gksUOZQXBN3mDTZxLs8COdBCsg//TWS5
2rO+93wyJOUjapIFwzJuKEN8Zw3UDsDh1cSyR0JVMv2beITknyZcZxkMaGZ9Sn2BERFbLfrhV7Re
plM3dzuXfZ8M9MGTh49ji1w46Uwm3uH9OWZl1997RKP7AO8krszWoalErzyovgz2VnroOZYMBVME
YBqK71ro0BxUMV7CQ/mFNwIUBZvfXZGzOCYelNZTi9f4FDpnYhHHyRbt79I/tc1G1tieDfN+03lh
hZhh8KnSoT7c4RccawECmmgBBh5OdjdROtbYsZoH2EeJIqpO/nxx4C9bMeRkXbgi/owEntiRuqZV
XJos7Dz/8+ZB0PyQTa+qOluHLU9cIGjaFy/uM6+kIB/SPuxmG7MPItN3mFUAGoRYnHiH/tYb0ICI
djR3F6Kre5/U5bVijIGuq6iMlI7Tc/Gao9CN5+N1BctE6uqYsRou0G0as4SBk+yqiV627DcX+h5r
R8EIqobf/gBFVaNcKeCIkKTM0j/qru+Ldiu13URJYOrKH7NqxqkiQC8omDwMus/UfbaA7t5J+8WK
FXzPxdV5fsu8uVEi96wWeYyxR2s2OdnLz6LI9twfsq0VWJ8XJHGVNkJ3T3H7euhbQn9d0Rf8eZWz
E0gL1+rnNSpgXUTRWWhyeG1vAoY6m62a54fizggktYb+q545/sOBrIwqIpkntfTRxBMqGrM8C2wx
M7ku4aQuqchFFFMG8MgazhSlTWjByq7kfHRXEBlhUGKlGxhty0iHcg1bQOg9kAuGyfF9ahyxR0RF
4xLDTTtJFv0g+ReLmJfm4HB5D5ei8Uq9fBJTRzJSc05rZyqDtmy6wBOSmPphV/CpABOAIrwHNW+o
3haYa2SbIFkRHkKEg825RT9rWYRjYd58liQJdoTCrn35nDAPtwRtjkaEtK7hYXN0A0ZQCqJLorB7
dBtOgHsTlyyS42CiGmBgMBoeqQyaKVnlV4/IwlyM2ciCxfxChsAUGLCOXtxmL9X6leg6Jgtj7tb8
UT9Za7rG+2eTaUOg/0gf/hYvjhChVwoLQkjyxoe71ONXz5TONWb28FR2quEOSSk7OhUaJIXBVvKQ
/FvgciEn1rLKms3Mfj6SnhYYojToDcSY4O2ewX5ev5JLW3VA8M/IRgsAjne3WkBDUK5kj9h8wu9k
EYgGvKIivdGLqKiekrzp3Os8OwCdEhjGpHb5cUCcmt49FZsBg5UL4uiMS9U09gS5TZDXqVEB1Zv4
hsAElcsZKH/byy1PAmZ29ELEyuw6oRhcQGqYBZKLvkMW5TWThgBUztFQZ2eVLzOsZ6kib7ynEx8L
n8tzzxyaXqap7oskjB1TK0nhS3jysGn0KLSsAH9fMlqDCQsSdQ7lym8dJmpOJl4CckC44KtrB8ao
x/gfLDauFBPmezd0q0bmmAN6mgtQhA8jKQb57nr97So7xotCIBagPiA/lLW7M46esJE3m9kE79BU
31H9XTuELrnTGcJTsktGuaMigphIEDlYAVEB2L17fUCWk2Q9VosE01zARiGJLcfuc30mfS/rLT3D
999BmGzz9MhbICMe3hCMMLkmGI6MKrgHC7ScADDAnGhkJrywO07GZrQ7a2cGcZfIp/yr1IoHwHoP
es3bFp7yKa0lLzUcliAyDX1nUhkxgnXuOmv5Seg48wwYF5dTuYHlvnHT63OtN6Uyv9Ye9QtkeLUE
6siDvOIVrgOIT1fU48nTzE3Ebq3dsQ6jIHBtwCHpAd/kZW+B1l9ysfmmWVks8dSR8WpyzzBFIwFD
SR6il8iOLnWkzWyr/4vqOlR7L3ty31dxbj9PpQVXsYNU6CbWqBO++JZ5KxY3bfThsx7Koof2A7b0
WrXCz/Iyc1DEtm5RoHxB/WcT08ug6D6U2r6ctCw/wYcyHUjVHTql7PyDdlnanDLDBi5HmG3P98RB
UqUFKA9+F4VFnooWI1WnD5CHO80uZxONQrFAfJOzYC4A/7Pmb29QM5wGlDrzDy8FF+NQ4rnfWM8W
MAtC8kYeHOUObdjM7hq+ZTkqwsvY9wAhzzhwgmbNps5DZRBhdx9dGuIJ7PGJyBW45jYpuNvHbeMi
ocadN+VIG8iIc+IpGH2FVcri2yOUaijm0GSMKhmC9NayV6l15dGHhvDIOBkQU9WrMQtYxHinnb5C
tljP58JfeCL+tf5hJNaGNPF54mknSHkyoGg4Jp5SmyrEanmfD315UczRq586nJ2IdEKE2wlQgyFe
0a+6iw0MeC156izqRmg/+GYb52tFUZDAIGSp/pucp5ZlusYVeqrj2T7XznKqSCcoFId5P9v20QHI
hA6aZzAv4SyuvEy4/UFAP2FJ4FFsMlUE8o4t4EMknHO1uCplh0xPLl2vDLU5pRcXsdGOYT33k4DD
wZSP2O3bCWkDpHYBFpwauC2Y1wUE9ZZMb8KObBMA9c1d35Bas+7pdoyjnWjVYsAJNbWh96n1jRY9
W9ZTQ9IEfHSVVV1A05n5yvwKilJLYefr8q42pgjeANUSSpx5OyL5Ws2gSdo4EOqFiCRY8LckjbE+
mIZFyo/oWyRAB8SBjDvDusfmJyQS0NKzCnYPi9PTquRNYuwP3MABitiLjGvPuj4iaoVlrARvAbGn
sZyYCioJF1VCZt4Yt0eNAX0D0rBkb9p3NwGWeNYSPSBNJXa3amy4PahgUv438ByFuVNRsPmz7VYA
udL6O4YRkBfJSm+JcuNA86G8ATyatLMoihIr5tc/sPY+IKKkg8D18LsJ0WrDaq6HfKWbKPe4ECPe
k8VhDM/msAsfKxPdPsZTBkeZLHKdcVZ6+uzQu7h91mCcMBohw8vEBOj31NUA2rh+9M1mlCvDTiTx
r6QI4nVg8BJ0Qk/8mvjP3WA4rmfyXy8+c3jHkIae2J4MZrQB8XMk9c+WaVMQyeIlhgX2D64zJsZu
mWS+rdmdkmsiUyk8RWn9OSejbTqAMv3AZBEceghZ/Xp4dAdK7pX5wXoAu8TGEUCd0lKtrR4pNIYp
zsVoTEzYHY8ZyvSiaqBowXbLriCCOAE3uEPdOIPUumQMHkGlIIFxSmMG4kZpZSZKSivhNHEZAuhN
TJWcAkeE9EJTeB4+km0k9JM306uhCYziT41dUexxMb7ub/ZL+92g/cdL7bTXcojjJ3ho2CrxplNU
ovLIB3aJpnHAWXdU8VJMJIOwgBiVzgfH5u8q3IJ3ZA2JRT3oTLnF5oWOFHyJhX9qa9MdV6YsB4PY
emy8bu3P7VIh3FiJsqp0yuylQqGpyFkMzLURLF2pW2XVJbp21Qk5YVlLkqVKizm8rDfPqwX2et8v
h373wnC1OhrVKmvc/Ju64HNRIiDO1usIQJgV6bPtNgSPmxKmAc8EzxrN7WK4gP8QAX9LPoUBkcPR
H90Ch+lw1f+URJPh+vU+5X6jnv6wmugrEYiYjxhwKaY36MVJtHlTgDP48Pk9uas7IOImfckxpNM1
Ovx4sJOtcDhVcJ92C1ExFKEaaUypWwcV8kzFJR9rARRf/41dmIXISIaZ45f8/drSqt99Db8TJfMx
Sws8FCLogtEVeHSbkzbGDsRaYN1CSRltaFqMY5mj2NGO1YCwidaAEKQsQOOI5zvTxYDmTLDC5u4I
Hwh0iJr+Twe/xYelbQZRQQ49x+Hn+T7QfEed5qDc9KdA+cy2890C4CQDhmGUbJPg3JNROgTa3Vg7
BNACDrGwoL9J5r6xbbQJK+xZ7z+YW/6ZVqMg9HUVf7isWIBXr6KddY45Jvke19drQvN8PLtm3BgJ
oGeH49nnkcjIMLh7JYIuDwsqKl8Zgb4FSEfT+agEfZx42l08vKpUWpjz47lMtI0sN/WO2S7fMM0A
3BhiScIhGV42ofgTA/IzQchm4FOGpfa4wpDBHxngBkfDAqH98EZEXWKGZOr5rZ22rVuW89TaEShB
dNmKuuKJ9dJ1R8hvkP1k9RCgxbXfI1JKqxvnWVBNElOT967LJH7obsve/tkf9vumU/C87XJKcjUw
YArcV3oPforno2HKrq8OGc2bz6Lh/Jv8OmBDFQD+O9+HnDfLJRTHlaTy0WHLQBfS07YW/JA5nfgX
J3LAacFCCyRSZ8mTWFwKYTnu2qeToAyqsYfBD2AfJvENcGaBQ2ewIFzG+scAcAqoxYaCxlzxsLlc
WTKURt2v3z+iSOBNrYiahB8SyLvzYbSuNKkPks/LTrmCkc1WyCeMWcD7IeqAetmMBvOndokR9RmG
j9gg/uI+dasM9EVYQhgRx4xYWVYVfmbQ1Dho7rCId94i73sOggunsgIYHA7UyLFhFIzapVHA3wAZ
4hzHz0q4J+OO7qi1B+B4U8wmlSQdv5ata4guAaG6rJyRpjHUt/58pLE8vYntg5adCYVGnRXOl5FY
hlFb6JFtL/Cgtcbe/8W480h5zoSC4Xs8Epzyez2XZrNJIMt0CGtd9dQyxOKEKV3YoyW1nps8ccKM
cOLk4n4dHgyxuoijxzH0Zpa93v5AYzKZIq470Dmij7Kb5vbB5olA33UvO8cxHuFb/6uzq5tLoPSv
l/fRPi5y9U1LXIaB2ajY+iEJ/9Mx8kNogWGIgHV2dQ7DXrKiDjPDWw2qIRAd5Np6PyiO6fahxXvJ
Y0t1QRFNsrvwdWN3nDR1hPdpAXdCji3yqIdVR+6NjYezWT1bu7uo7o4e7NOSQaX4p+xoOnwXNajt
5QxwxrC2zuLt1Vx5HLlDsaO4mBvwsS/tbYy14daV/ytwXMWfUIhUja9dhvc03xQjhlyR3Yn9a/Ng
JQj78xCD5hqPfjbdn5kgB1wNhkpfTHB3BM8sf00JpS8Vc6H97fQuERX9Wy9Ii5AK2mAS30MaVJq+
ECtwC9+TPvg3S5Z8uBGGvuoV/iXIMoDMxXBGgMNcTxWlEP0TgLrfnwOWa1D3jz0dfVj9bZXHAfX7
DP9HDP3dA74Jhb9+HlarRews8VlEViSsBS1RL4HJrGxWBoQ1/vKgHCEkQdCj1+M8QBgRIFX6fUyX
NvLEU55rrwpCtkwVb9u0Wx9H3euvahEekdL2RWG3WypQ2/ZxFvFkKcR81h0I85ylYjlgxPcwizlX
EL0L8jhxu2NKS5E/ea4RaNgTx5ctcnp+uuvqHB0vCGe2nGO2WCSqTj7Fi3AzmhsoWJxhpDAmhHM1
OsLHvfeNvwzyg2PVukO3J5f8XvgIyNi0gbds7cU3usYduwTipTlon8oApbMWkjiXJCSM+kBvrxTS
v1ark/Rg1G5xlkqMdhKwxaL8OWidp5b6FFMdYdmqEr0GVfmNtw0eAu4RV2+vJ3RvTjZnc4XrKO4t
gkppsxj/4fC2tHHQh/vTDr3H9Fa5UnbOd24AYYX24DiQCeRAKendFNC1K+Nr4jSGfHXYL6K95Lgl
+jRsPkvbQ4+eoyG0zXzVXNxhOf5os3IPlyjCdpN4XN2jtbhVaTBg8/kxRV3sf1eEeKzYtqGCcdYC
cdSZDyBb5xYh5FQ2T8xGRaOzMUbgSTPJS3c1oQckwUZQVw3oWSXI/1aouSZmiN3KA+XS+mY080lC
9FGbgvcXUagLZj3fNyTf7NIP3ILWTPvk/ms046BDUpJRLwt8A8PxNQtUGBGYCRS7PLHRqXqeF5+d
C7ZL0v39BqBNbzjM85s3NY8V1uUqQ9CVIB+73O5/aVjWKDITUeHe8nfYMDqDspTtFbmMgsixnKay
CN7fvwrARioko1305RSPU2o2yEA2Ms1uiaUFWu9cJJo0jA+wXfC6gVz+/EklpqbOj1UTseMmwi3I
MVDuT7fdJXxXF1X3VLqInOZVWv0VviOjCILj9w0Jpj8XQA/P4zUNHHoraP2HsL9UOXl5g0lTB+OZ
xc0nrlbGEenxfx6ZdiU1krpQ1MeGQy+pY2TcX3n3xeTxZfMkHhAzSZ4Bi56Zro3j6WhBd/H5GlP1
hW7Hd8HTQGO+/ANoUiHDhEBoZqkoDH+N7dZGSDrCElASXKBGBAk4W2KoFRIbidquYGctRyOgGRCZ
C6j+Pem9eOU8pyD075x1vESX7uP9Oaw67BcpWpVoQ6mnJnEY/wHRxRuf7DhY6Xsk5rMi9tdFKhBM
NmYCbgZ5rkKSkF5j5E0DMsAstWVQYnptnvDf1/Zo/SG2VwCdX6/BmQeSwNAnSsb9BWCd3+XYTbw8
3bFd8ep16iypBMeD8KWSpBSt1QD6sCLEni23pcSjDvhwHNEmLbbI2HFgvx/nbQQBsrOqwhB63eBb
926ZcAMcJgdkCi9urf67PQSaZkgWJDz8Pa55JF9xZdPFhFyMaM+8ka7NHmxKhtDC75Z5mm470SzS
1OTsNi5+FvMqjDBDyj5YlorsM6LZ7oIRl830F/kvYS1z9OU8NO6HN0nfm8EPTbfnxSEgO+2vXNMi
GoNEEvD15g8J287arDPqLe9VBhHtMn8uBOGs7HFRkIm01yXv8+7OBaxANp/VD8k7P8dUUOjNdaLu
Le4oGe73Y70SLjizIRgTl2tIG0Ti00CZPSWEYDpM+N2QsAM9HlphdbHiR5B+s/3ufbp+yLHqYsuS
wB5OMMRMlf4VC838u+9p4fqjUYNPAjDEVyK2iuOP2zqkaGygFvTkqeqGUpVuXTgAXfpvy74ayx5p
l0qBZ8vwLhqvz6Bv9iAJRKLIfGLflZBtI+eixviqkuY/THuPTjP5xOpx4wog93iP+3M0KCBa88f6
kD8x444gCCIetaHVtb8n9KSkX3+PPDyCeiN0HjpbtfmwsbOcfPoPhyXR/AwkLDodDzT5zrRHgfvo
IbWqA9F9TCoTGbN0biaVpei1Nne156PA5/SKlfOLMX4+LPqlhlKbiTP66sZR4fjIWQ3NFjdK8Drk
PzDi9xyISHzxGZjhmHama+79v6QU9WzQPmL5osjsFHUFmiJn+STb/++v7N/pNDb1vY5vh4qZylO9
rbBQQkeute2U4cQzYtreE0+alEXyUHLYOlIfKzfHFyhnB+/5h0ZwHbs8ii8Y96lzZCU/OSlThh7S
s4P0MwlnnXz/8thedp/LtyHp6/NxaFs/VtBfHI7keuSbdLWWWrKkDVscLwEOFM8OQOmau/zqnw0X
R6/72g8FI+jhNbTxXprF2wla/s05Gnn6Qqdfl8qUmaZWfLR/WLUtciqK6cW3fvR8lTZKA7F0djXY
47Z6AxS94+/1eEyIpUcuL0Q6B00R/UsbwX/JEXr9ZsNIP42zw8WLgQnzQStojDBecZIeqMnoGiWd
q4aYvP5S2FccGtyZk9EkB6qzZnIc9EWyrx+OX5WYLGfCroCFHoj3LhE96iRBvusn5cPf/uabLtKz
x9T33paXk2HpgDzdbiBCVoLi0AtSR27CJYVGD2q8BEbkNOsi5CpbVA5bWq/0mrqYTJot+JB2oZgq
DNBi6m+C3fWu/ZadvdCxUEhnRhpSlRt9vIhEIUaNf+dFhfyxTfy76ghywUd+4qvkNC2DdSqnBnfC
AUNmwR+i7lCKKugYRS1ZFApZLevf961IARfqo5qYoSKlBFtwMBnIv0wuyW9ZW28bXbvD2yXivnL8
+QWwrF1FQ9dpLwgeKwRh6jGXduU9pPXZTtiC4IGqdibL9eBREdzxt5rXmE8Okb4Nciicd4OxYjDP
kf+rUOCrtyD1aWR9RReqJNObm0siK43V/nwCrGaTkMlcG3/DUQUndQylud27ZiRg6xy95+EuMQkF
hiaV2tkTskYGgwj0pddbTcAxLHuSs9hvVDNIWKkAAxUd7iLO6mDaQ0TbYu35hYpAjAU772oRHEXk
323AKKYAzW/vflKaPksJn1tA0A9bsMXijJivWXSx+BMj7CqjWhIxzT7wyIB5TyTlOfm7RbWGwM5W
UZ0JDdJT4uxEFHuY9b6XBUD+0h47Eu6xZxkq6n4pA0h607UZ+bp6rU6cIFHd5IqItDm9rgvF0Rc3
s/hviYhDWh4JmJwKh4xKtbL9nxvTpfMxVSzdLgfg7V9mnE5fbfkFPT54yyPAiBSfM+vjTvrkIE5i
D6DSkbJiZ5CByKBoU+Y6Fa5ipADVFVID63xRrOkuHBiYwuRN9S4B/2y1f9k1hvetAl4PCHvGxEQK
h4W1MZWCg22urDIw9ctYLeXy4jLiZa+ShCNQZT0E/zwhyPgDH1nfK7qCPy6gP+lMbDPAXBlbvq6z
wuoSPUL4UnsEzFyVwxIqcyaspPQqJp/GDeyvjPOEr2nRNfxqi7jaB4AgHwVDP4nJwSbCxN5DS5pb
Vj28xZXk9qXFOwC78tYxroV2Xks3hjurFUhM0fyO64Bud5pyO2YONDTslhGFneifjKBSsgNCqD2M
YcaRyuZ8Q8mkSYnYS7C4YJ25lmAdflGVPaeEszXcy1jep7KzMYD/mUFJLzOsTarxCwV32yNUlS17
lM+dRAPheFhW5k16mmiyNUFcq7di4slqcAFLOo0GcoY1jT8rEbabHEp1n5nbld1CXaAB81CF8SbN
go/Ov4KPyR1OjZkb9xu9UQR6Tp6l7XaR1nZdQKwiX5DB6hIzRagX8MAvvxg7Bx58Ja3o20xN8/uK
eW80MVQ6odjKGiSs4ViAhZVeTUIrSGV5wCDqO9G8jw2czYqUtothT66crGnNAQl6Cn6UH7Jtt458
/SriOauzoXrocUApfV0qNjXPe+dutVjgX/6BUvqOb/mGVyTNzJQXWrzjlNaYgrHwExnoqhkVJpDJ
pYRZpjCgrfv0ZzgAmteqHlDI7UzmYE2SlkJysPLYjdkK7wcY+rT3rfiZowqqjmhRZCI0GAn6uLZ4
QLtv19Vr69LwGuxHe7e4SqEPXWE9r++/i+jVZ++V2ZHbM1StUcGCUOmdm32JKd/wIINr03PYmfFk
nWj1Lxjtmhpvjlxi1O+deNILgU44jLOsJfIY9kdoNBzYowROfPCWbnXrVwrNn20aZv2JVrHWNlKW
sXpTKDkW6erw5419rm0AwHBj8U0y+K0IZ0Hwt4hZiD6mWhVbScvDUe+gu5c/Qqdhi4M7ar+TrFhT
I0u10hoc3Jz45evyTjiuqyXaWGo7MkXd/cusxiJ0p347Dq4Lv/05Bys2a0gCegpb5SFljqWiaFbZ
9eYdOyEYG5OQb5dmqfHwMLFEjoKtKcNbF0mREBM0iMRsoVBUrKyDwT/KUl4qV92TaxQZIfvVkmDA
J6N3gcTv1zd/iiPYqahxc7/rojDkXvH8zGdS7W6x9Bl7pa26+UnZlJqF9TS54oI+XI+1nBY8iij8
Y1GNpLooTsIXcNfkPSZVVRPW56O2AyWEhSe1GuK1YtTVRXAZHDhReXn92g7vd2K84S6F8N0+C57t
7v9dt9Vb7Yi2RxGC9h76x47/jaQW5VrybK+T/E4GzWcrDO8+uxr6JVnhkO7QRxrXWIoJ4Ef0fX9l
JEYbfQS1mCFmW3fviPHBkvMlDelMgQnXuzSFPQ0ZMaLDR7K7qGJWFDL3+kWxkgKxTrbT1qcUjqw4
hAYAbqyafewMptRv8CzSRDF70b6mxG1lvd0i86WddboGuyTAKMPLvUKp2FpdqWt3C2EgVmTISC7t
YBaiCmH4q4OJdNjpRGQIfK92R2SDUJ+sk461jfz271DNPWQ48F8mQ1hWSh/nmCL2Ass0K7AT4RNF
ofcrE2x4mcuQ4DESynpOr9LpOauVfJI59oCJPUDfnaGgYOfw52COTuGE+StZZeZVOG2Tk/sYrhdZ
DjTodM9dVVTajuejLYhXeYmPjw9n3q1cYtOIYnBiVTuEaxhycqHJacVeHviYZp0GTikjPWOtt/i4
Hmj11MHSCWw0KtcUX0lyjLox9m9d7+7R6qLwcqEsjIjdEjP43nVBFu9Ccp9qlHb+VThpQqkrq7Hm
NVqAKli69UnGNNwxm0qrGeKGNrgGEOSN8VfEMs3nFZpsXbKtazuTblTqNGlx1i+oc51TWA3KySB7
fXT8htf7Y9yYV89IGgRoihX0bVBjHdWxvNV5HDC41SiL549/AxktqJRYMtAYvKcL6aMFLghQv6aw
QtA7twztk9pp1dYqQbs5gzSYBCPjhWtcBdAkUmvnjAGrl9g4ta31ShHi5oE8fA4EXsUhpKn4NN1T
9n1aObhqCn/rLcf6IURBZCbCgCUYD5oroiJ2MNZuyU4Pt+pO+Fi0uUhyfDCSkEKvD/JuWv3vDaQa
9LrIuS5f9vJZalF8CIYgIENYKgWE9yKO5YMe3CM1Bfn4PmbAUqC4XphOWmKVxUCGFYTaFokwKSz9
b058t1TgfYFBDCCxdtgoZJUGn787TytU42IlCrM0+tRH6fnX0joC/3EyVtRTy4gAsV54vYzooy+g
jdZTTqm07k9XDDH21LNWncwo+wGONS+ZIkdtKXm/G6zjaEEDA+DRgKD0APqptfE1fOwwKzOcdgXf
uxRdpX5Y0KlOzAkyEDf7GNpeKOxeszcIyuHinIV8zROiH5TsE/yGLUABuyQwI6Z54kgjUBlla3Bw
17PZukJYT9fpIBbLMBl1SemZpbgW6oZ+Mkht7ghLozu+EfkHZDkepn+fbaKmqEYF54r6Ii+/lkbZ
nf6UZlG0w6H5gq2qYM7yGwbv7A4a2wlcGyr3j4tjjmFpuWBHnN7PngAESRWeO12NYZ8OpHIeF/UY
AgWoZfl/aVPhhRnO9K2LQsLHlVlNXbheUWJNsUWM1jsnDyvUNlk6oJU0bZ4WuXhViXhGm1MN3yi4
NiaM2CEEU5ZEolMQqe2uOJPmRiH0mEoHK/HkqaIJmbHa/D8dusxxik/77HAP+kZaO8Em0bPKNSXC
8Bu76Y1R4p/BE/xjVgmWnCi6uzzkj/KGNWnYwn3YvwJ0rRI3ofFPqe224GX6YHoblrRAnIh/CBcX
gg/rrpu4zk4jsc1nm4bN7IPaGy3FHSqoOhx2tcTZmBZk/mJcCbEs86bhZVbKodbpokaYZ792IW5r
pKTW87PI77wifPd3G/drraURieZ/vcrrU5q45RZH1w5l09i0eGz4g01ELe/vEbppbv1d4194Oqb8
cLj8+F0ETEgyaJ9l0h2HNkMS8VfcUO38GJK3m8rnENYmf2687nfmMKTo3KRqlh7hDDc/TEE0F/eT
LCAsxic8kSm4yUIWncppYsFwvq3hJR7up/kRvkmIvohHDN7jDoeGnS8d4D4FZAZah4U7dprmdhep
bIp/RXY2O9ZHc+DR7WhM1XJlb0NZAD6jRLEANvDcimuZ9ZrROA+m8ZCWxvn1qexbsuxriq3b7w5E
vC2194MyHp2H0V82uCSsW3K3Ej2MpqzDSnM0VVutIZNr7DLhvO0Nr2t6vFz4brmQ2NmHhqpxl6Qx
CVHTJRAVFl9DupJwjRYRblPQSlUrY8jUHy3kWeKdKNBA2Yp0d4QOb6LZA7sD9RsnDDjpvUF01Kjx
vtIo6brxjwHYIl6TS8EiPeDQcD4LdeJHHN2yDFl2nB49czFYsMztL5rfUEryoALBEY1dBmXGpCil
svmajz17Y3bnYOB806MEOom88jS6rPpHH77yOB6gfm7JHGjbK0fldaxubvRi2fQPZ+zPqJvXwVgZ
sUy0T6v5UW5EZjPFG+zdprVNCQXNj2e9u0Qsra0lx9J2dBSSMdKO6VzXzVUo07ljuisRvfXxTKH+
Z1eZTM02w0r+dbECA2aHILHZpovJ4CB+QhwC1hMuSCJlQexzHsPNmiRtS5K9aDZCQcQ039dlHv38
P8PbfoFqt6m4yvG6zYw4dW1JnTmktnLtjjRM35EMtqd7Z5DdM/c8Ce7n1gnd2eQDCqx3iVSOMVvt
Y8P5rRcpvEsfYzOO0fkIKOaloVY4MF+PXzUr8PrOn7GC3hD/31zKspzW8tH2YdDCRCR7BM9T5lUz
lZ4W9XZYKcUfK29aIHBxzZJ45Vg6fzkeV0FjGnBVRokkF/BHdYIZG5nwvCmgGNKOx76b7fK/+aYz
b+50cDoKaYTmrs0/lR/yIUThBVy2Ev8FbxEgxI1yFGiGoC2p7VOTgpwZGdHedj1MYLVw8AMDcxOP
jFc9hJNhg+KYGh+lqNRMKKFEoKSTDcdh0WjiMD4hkGXqj6zx6m2QpNQxwbXw25NjR8sX2tUE+tQP
qDtiQPRsjoPT7GvXpOkfArPc1OhEXjW8w8XsfYBsfRlvWYZlALPjg3N0ZLpIrPzcHkWHWcFfn13a
UASEi/2FrrpUo0ZWBbynhv3xGL0ZfB8z3NwkG0MQrTqPHI6wAQXZs477Wv3C8Xm6sVexZCk2UA4M
TRvLjgaXsYqd2kJtdzNrXqO0O63yPxWlzJB+ZIX/NVr2NE1gFqYoUQA1oM06urrObHudXDbUQdDI
Z5zFXCrb+Un56gkX0LuCPYVo9YMFS8kBJK73y77lrPpqTNpf/71oS500765RZEj/asp59n2NI3QJ
xJ/fIBPXT4n1zK/9wLC3YKshZ9/Bvo3mknZEO6ToM+0lefDT2IqL+IDPzE4VIAq8PWi3OcIVxMkv
yuGf0AJFYCzxOxhCLxc5/B9n8KnnnCKqTwckxdtrr0t+59jlzCWbUuD18SER3QaeoDyBHKgdBJ7Z
2CokZn17+8zEVAmYcVrhaiilkA221AiaWZMn+wSWJaA5aSCIsozwDgn+qW+070vNjxDgNGHdnJ07
aLG9S0lUeNmKUoQobECQBasOv6RLRoV2SZSXY9kxZspzLQzV8u3NrBXntqWUa2kqI8dNv6UkmXpn
LCvaXy/ITYHSVZpa8Kzpft/cM+7sv6hgYvYCXI/WSZLzHhC3uFhEj5K0K8InznwquexFtXPl0iMS
Dn6/A0e9x1r9TdlRqIDczvnFC07OdDq3pz1AOWK/ZRza4WuSLZPLJOa34VbZ7T69rsTS978rampY
S/l2fdLQbDjGB4rGUEHb3WxNl183IPU9j9gqsG8rp8uRYOILJzyFd/JmCzx6f0QR/y7tH2pIXlI8
gPfu7XbKdTADLoht3f6Ioqfi1tF7O9if568jzS2QvsglJEbqOwH9HBDu2VP3pwiOECeXRJMZMHyq
uzH4uwnH6OafKzclCcuZxZBnJJodizOB+WcHpoGfvdKdylQAKNZij+wRpZ3yVMRFMqoa8mxnIQKt
4blB8/Rcc6qh4C+Mgq9mjWAZGtdcOnxfJLDWG+/tpIseFQgokqw0+Iu4DkIqQgJ4z2W1Ns7GvNoD
P9Y583+B+vXLVQk2b4+wUPlxRg+s4RRcQqjdQOZHuiT5o9ThHZa4xUmXL78QiesKcktSQWXI3nTc
lPsTsqnV5tR3Cv7hEKrV8eJoxKxoV8fqksZ6A6+Ffzbk+EHxQcUB8Gh/j8hfaYJDsSPusSbp/ELa
eI2UWaV/jF+NWdqkw3NDTh1rgpndxfXWMG1SGFHyrYapSrNlUGUw5TWLQ50YKnqh2Sh2aptN3IOy
3Pvf2u/lzANAoOURGNsceBhAsSfUZZxj2YZXWMSfKqTr0TGIqeBEnAjWcA0yiG5/xesu1lv70/U/
7V3BUScRUcfv4rtqMiL5q2pGOrPTt3v0sD2SiXYhHX0QK3ptxwY9mlyqHhD4GqbqgAcCXWhhNuVV
anD9Q541ps89rXf86lhmDrErzIXVXLN86HWTDJHi6VzcOojG40ikeyNQ0DQPRNboSMxj2/fGJxhf
eOKgYT/9ckymhblSlk2D7q8Fe5UlkA4SlmNPzv7hYCKPZtmd4SPIFw0pavJlRXOnRE6e6eTfSIvq
lsVOlOVlDGQ8ueegGEKBWLb3tZYMpjwFE0XxKwHLhISfdMmIQrN5sHGMTc+CvswhDkVdKau/kEqI
NK5sIJPNLZqWusM6deK6r9oHvAfqFxTHAfl7rTauNADhJ6VNSJ5HdYBkmUmFyOvHjkjtIEdefCf7
Mf1DrP/44oGmx0stHwnVGV+cEkWGq6ETbSN9KGSrySNb0um44aEuG3wnCxKH9+CmgfftJDOvWllK
UfdkfmLsVH7vHlgQapChhUn708lzUwUvTe6eBhktspsGS3BQ8d0o90y0YKcbCFeJ/shgkkmTmRcl
n2+MGJ3iHdyCo8H2Vw2EBwuN8W/o85KlK//bqRm8bOeyAFt06tURN1IyeerlE3UeaToAr1aJAdnZ
tawyNWQrYQ6QNbrdW5vOC1Cj4+McTWsKzFhTbkCIPBfB30Pscy2GcUQ1fsEzyeWbhLujf8Z9/Tpe
D/rqhx+r97uWM5PMNOMOdOnKeiICC8YOJRS5nfU2KJZLqFi60ev3r2j8uE74KRBSw2+lEhic7I0E
pU1VEYQ3MwDIzKpjtJsuM2uf6HLFnUvfYxuQyG1BiDLYQpSrZ8/7huR3jE2mZpYU1U7IYw6ttPoR
I0YO6fLdSgjLIUmMF8kpXKBx7UcjAz/1VrLQ79zxWbvhwPEXkwjVNr1YadfcU/iXu/E2cJOnsc7K
lU2x+M0KflmZK7YUmbAo0KNVABsKaaWsZsPyfMFbYxxOzr+ESojxTQ+dIx4mGmRAHKfvE2I6XuRw
I9L61ZcO/6HiLv3gKgM/nxiLoHZFZn4Q41evGe54kee6/NOSkQxJ0stTv5f/iOiBbvnrd+c2Z7pn
/gaey9RAxdsobwR1q/zB1V0Tz9BtX126JGv5T5MYKlKD7bI1Werc8S3P7vgYfxAb5uGqCu8ONlbl
GhH6fMrfmlrz0IcqtjPzcztYN3gY5l77GCUy9UNWJngb6VS8l3Ax3ZVZ8UYFBKhb7Igl+5IxzHY1
prZq0TO/b/XPOSCEMRH7B5Ef+h8IOOPXSjk4eKpS61dEI/yXOfZj1acjE0Y0QeeXZZJ/fWf04Xis
VGjgxOzDKBSz0DXrVns4Ewpp+5sv/33WLA/FhONhDKBAy6WqENZaOBOj1mG/rsTY8NYFIGyNPfmp
VKHnIeSgrf6QKLPGYSQGEFxamDP+vVrJrf/i/yRhUHs7wpCeml5yBVz9xGqTsS2nHdY98Wm6XzGc
P0UWtxc5VY4BIoM/SHN58tQ/03MJiK0cEpeC0hnv5+XsF/GNGxqD3tEzgqswyiAScmIJSGGFiAiS
ENXd/pLe1/+JwhVMlmckBznzxD1Awv5LHDJcx4JV6epTwS0AXVRG9s6O7bPqo6ltahzsIVvYttVN
1zbJ/GKTffNiSFbVCnW9lxYkyRAFBXfFUpf2qOgjQIsX+1wOksxcuJtFF162uDYqT50fv1w9gE9S
WJsd/zDsCh3ZfnjMBN/lnhouVKsANLtu3Wdn93QjGGLOdlgQaPYlySUAPBWh1TS6mCOBfKMepOdY
CdRVb9XCmjW0SqKLi1NFYzqAupSJEc7AEdy19afSUxaVWz3gESeLHWuYEU9wuW4duCsMdrrSHicl
Y+y9h5JS1Iuh2LY39ThYWblHmIqjxJJiBNkcjmRmbGDhl32eZwNp+QNRWlyiwwEF8BaOFhd3R7T3
g3Dydkbe6zvlrhQqRSklNUY6Yb+wJBtsLGI4KY46eDdZBkUr0eJNIby33Z6gJb2Ym7lbV3Ivhhqr
ExgYVjmNazjNbjmCFCiq6uchfWM9aTH7ukeEMHMPE19NED4i9K7fs+YFCtHlAL64UAhfToDA/8fj
W7Od+vpkMYh9pln5hJ1lpf3ZZ8UkkYeSDzo2ygOQtCxI2H1+5Swm+yheXJ3EwfdKBvTy6++QLZzS
0b4PpGj2AkgKd8Rg1jl5LASNVlX6/kpPiULLrMnx6ZtkGIlueUzLGbU+kX6tvOeOmFpPHxORw/U1
iTKS5ItUgfWyJ4IJPrqWjZAMvTjS4SHapNdGXrjVX717dkWgpYk3FeDyXNwdPCGlUPP8rnjg8PLe
ZRagH28xV81MWADtKyZtkEfFzMWL+KhXb0HSSsF1s8H74oyi7E4+Hlw52gf4z2E8Rw98zGydeYBF
una2uG/28WHNc9W6VXX10j7iLIwNjP/sMtG9pUnhF8vlMrJMwGqpzLqn2GC8jXH1nMwPvsyjvzXh
WoaomTp8KX7Z6iCnrT75jJeWFoyoW1U8cXZdVKdBiQVrBr3Ph6RB6tftfS3SbedecttZZ9H0Xna3
UATGeM42LEpbe6UOZEs3Ge3TPyJOijIKRlyQStpgulMCVwftjIB5LDH70WUYAX7JrdlwYnmirh4h
tv5wMuXlVp/oKqddfOu0BK33KB62KFao5HGw0pHDhmn5An70CRcSDNdFVddoeKMtk/kTDITIahu1
ygZDU60i1vLZJiHeQo7U84rEDmiZNjC0TZyuPNFBKGN2eMyU5flqRmLMCerTTn5ImdfJGOHHHh8j
HhuiGtleaFULC3Ohz4rvFdeQ0kYL31rN674YJ+de2BXSaD3vehlCmtGistkAcMl8PWY2SRcgTauR
5RCdCgTf+3RMukqkzhveD+z6Kjr/KSr20lb0Prh4QmfYEQzTWatf3rJBa5sVrsPxeaspFjG+B4qO
Eejvr+7Er8H/198rTjU+5TZp9BrCZzegmQ9ppRQUmhU0aqCt5gqMrgIX6vp3DoE700sgg/qNRUVF
Z9GrgGM3SxjVdFEkJA5qBvs0BBynxjJbC/RjQBoYB3vxXe+7T+qIeGmwW7GcjHqEYutEm/XnRCLg
2bPPibRaPxYz9IUvPUgPjf/F/TZzgpycdxeHo/nBCZhFNZyHW66s7vgrkUqbVrQOPImqTCpKG8mN
4EtFNgFqFL9VSwBGx4bFer6Vyh7Fk8+geI9ji0dI1BFnKl5Nz/1DqHTwsUJPnpqp9vuGWEcyWMXP
GdAr8fQQCIyo7J11on8CZjbN9/QCHHK0sMI2QZT8b875IwpZmHmQ0PIa7Le6AVWEPQFkc0KyOAri
FlgBWEBelRYotRaJil8qU9lN4fJYWQbdJN3UOJxjKEEOaSrUKN9gUhOUY1QepcLH8wLuvFvbNI8e
6R+xGIS7fcAVUFyiNiquU/BvU5Sk3ihz2Upyee6qJ/BqqPP/zSDiyed4UbhoaS3EjwfdEnpcrx72
madSecNl30wUY7xYhp+oczbl0mdVcpIq5PCZ2IXWIs5qMuODFn8EPQGptH0yFUcnYqm0qxDrSmXI
QRSAu0dhBz/b0VV01aYC07XuzbmBUEthId8dmdf+2u7Sd8VxKeg8uTPcVqYCw4nczywUJ4sN5xGZ
G+KEpzz4ZsqT7AUh/u9MSTZw54mRkOvFsr+T/uIacT5AGxHVrjvTIyW3h5Hi8Y7l1WreeNQOQ3EF
IfSl4JVbCf1ZTINAM97Kh7aqddTx8KLk8GEU0FPQ5WLbJvWFpSAGlvCzi3fWi1FJ3jn8f+42Qm7I
C8uRjDvrLU0ruSncPcevRebl2rFDd+o5FQJexjlCm016kIlASXBu/8OC0+FC+bsUw2Nig6k2sVqf
9pTFAla6IC/Uwg4n7jzW9D6EpOHg5G8lVc0M3CniU0iUyqidWp3QgHm4PyHgfS/L/T6CyiqDITyF
0IPOx18K1VJ+oGW4Q2mvUxzrjIPrwN8YiDmp4wMR5ADppOVjmfMjkkCmPCwQAtTF5klF5lbeC1jN
fZGWqeZTNF90A2XsCx2rGTuhzqF2VBfcA2MoiDDYImjCCObT4GvWIGHi14T1xyoHQFaEafizO1OG
2mnAfb0/BVCriS5asGcGDtgqSFQzRsB7+NyT4chqjv2OfaBc4wYiiL3LLUc/SKOJPRO42rceEe05
MFPtTHwQGMH559C/M4KRyUGlTUFfcQf3Z8FxL6QE4LNByJC9l+gB0cOnmUAGMdm/qRfSXMf/38hB
vuYcJoWPSr0iB+pDK65ZqdSOhDprQWW64FU+Zgi+094Do/mt5w/c4ZNBQceFtGHOz2gEnDwEMzxE
rSzSs8nq8kAUTZAIx8cysOt91vAPcCDN0bSkHMXjLtZ1DxwALw8G1yxDRDYOCY+O34qxCxIrGCI8
GA6GOey5KOX46C6S7I6liJBUXGzIt7rrnMaIoSVoeTPHF6hSOTTcxEE5Ddj8fnHzVA53wFFgi7Se
PmBr5S1rLwSDeTesFb5KBn4Xq/ri0kPvVB4rk/ES30ZXU0vHswF6BJrC9Ir3NE2OduxzlDOCaYoE
UhtxF0R8bR2B4iGYbDsgPsnz36Q+EDNOOUmqnoVVb66ZqlBteogpGQe+8dhuE/K7+QH6aqwP97fT
r81e0ar3Im0AOdrC2AFYWKycwtNIkfZWkEKc49zjK8gR5FpkVPswzJorc4oqrkeco+X4RMARNzAV
MZA1wmPoJLnxZRHwdx3wz/u0UyvAjfJ1mauQY7YaEQmryM9b5qj55JzLoXS/Xje/jktPYm+Pc/iG
kBLxJ0BDGb3WqI7LW1fUC5Ka8XJBp5gVaDw4h5j2v9H6EcC/ap7ALHZaSz8CW6F5btMHmKC56RQb
mPI8nq1oUKBnFGsymiAqDQw1aBwDnR71mpUgmnJreSX7COmKUDmXuKDD+YJBqh9603KiDnWcIdHZ
TxACizyP76L5XAQtKgUHddf3SMkYs5+k5G16woC995Z/J6tmgBi9PKZq9ntaQ5hDNWh9MDH1uiJI
FrPLw1b9Jw9flQOzCREk/g9vMzbNyQOmNDqy+Vs8SeGcW44ii+EGCqVomHV5F5tIL3FpYDm5FVXl
5u2MFSUFPLWICjcd4gSqrk+XWLQRovxFCQ9zNIKruXantlTVlgL6+Sroc2cKSn5kWnSPWHMS7mCc
YgAbMi3D4nbQbbx5YGjlJnpN6ucgjMdAhBU/oaQjyvgMsE4uqOmzrimwLSDJ0PBF682HD6RD2EsV
FuX20x1TN+H1TVpk5yUG5byHu/vux0NovD6M8ZqzoyJWlDRBcesEm0L8JI8dQY14ssnMs3itJkPW
+AdGNeYvIdqGp/AkbveK41vKp49Kd/hwNPQHejGqjsJqmMYOAD3Jw2EVm7S+mIKnjpw5U+wYDM7v
jYo+DNPUkxONyPKa36t+dMq/iSnQoCCREx+Rmk7zd+80Aa+qoRlAU5m6i9QF5y/3AJKEulW+7L7K
tQvDxrplFzTkWxDUMqOAQinvgNWLuGXyzAEL3scsaCmFo8vZwhZ8kPYeYFezAMYaiDjekCBYQhul
tRh8gAet1rRJCKOE1cSoE63l3QTpgBTQexYVEwKmzu7YKXK7nZFxtpeTX4u/qsThma3DYSkVQ/cY
aUKyEVWj3FEFe8B/temAtFRFIUNb0PCxQOEDP/FDUuqcWOP9VOr40Tmb+OudEuOSndo/2AjGbJMG
mDfCZ+rnJx5zT2qmrbu4FRg+ClvXf9dX0Ppd+CIJX2+8kNUHdLna3J2xiRx9LiSQO/5s/syxVBRv
ymoSBJBbZs0jHjGv9gJAzORqUGtgI83TRld0sFSuKlEhvz1nWlCrWvgMFm1tHiD1T5+Wig8kS/KR
S+k87TcC4nz94mQPH2YhdPl6FTK6fZRVeEfTGXD8tfxGS+pQEJD0n5qNLdENNuW25QTqdkT3ifE8
35zFmP0dLh0697hhl+4oxGTOG72Jys5QuwwSWkFDPahqt52uj2dEdA4P7s+qnpPQ9Qqa6tyRL6tu
JZhoxD+YJjhzJNsWNzYl1l0UNw43sojJzZn6G7VG+zypsNA709MwnrzKlMtP4R4ob/6hDZOOliOa
NEKoQoEzGxS23fpWtkGEcPz6vbkPLUmdS3PJYLr6DXJ1HrOEEPqMEeGr9B5eqhPw7SqJhgbblZ4W
vgdNZqYnyBCgaQmN8wLCn1HqJaU4f5J/i5K0xb8n+u3RgAmGjZSy+Y8b5G/zbiMim7eHBQVkYUr6
laiuEbGdNkx5yKKxlL2GUwRP8yK9pvVlfUokL8D1u6D2WDGAa9FDXNITXSD3yqFQEvUSPuUchLLS
xPb2gYxCrgt7zvEoEqVSp86+rzlpkZufvTaDX7jNPJgjMw/gHbee203yYbL6FqqzeOxChyLKa27o
HiJD5si05zgk/D83jhA0J56p8cddBUNEAkUvFRVxH2na3CskJffLC3RWq97bHZbQUK1sbUDrIqTg
LkBwmTfDcZsdeMhZwNfmBMZVCLTyE4fFnyz07rloyCBS3p/1tMTP7or6g2Sqt+9nHoHOVIaXcQYP
TdxTC0YhIZ0Zw8nAp8oDmIYGhX7pleM5/bN65XKpXTOZt82XvPSe0gUadHYjfT9wFfYnT2GZkRie
zOEuwf32btO5H4IN+IxKNnqyhCAdDw0taz+IkFEojXi1++j8SKmLK5Q5cCfMpTZke19oyYwdcvt7
KMyHdbvhnlo/uzsU76krQGSMbeleQ0OMXV0ZGUlEeZzv/Tu+stk2LjgSTgX9r/ZrSqSRVRqcDIhV
2e2bx53qnCoshFTC00LpJQHAG3YJ4j+JlD/ctRGBq935QFI81SXEu+c8XfncSWoYGQI/fDqToROV
mmDr9a92iKarZjFMdCRxZo/CJ8DLM6RTMErJ8ZoUe6H6mq23ubxAb29LIc/6eRtrgRjDgIHKcb2g
J+YGNo5A/4ongCv1Mtxz+12SdAN3tNkSy2zTEDMJC8oTJvWLlvHGvD/0hMDCe1Kbfceqm7qMXAuP
yycOP34r60u9PpW6tedmO8nJspCJAnbFI4X0nOOZk8q8Q3WWENhZMEIN1dCKuRxcZaj6jTcZ5qc0
+Vu7YqghZ7Pf+F9k1ew/dPusnbtQnHNQL+z1pg0wNBfD7QPTvuPsObr8q0eX41Bnt7J0bx256UgX
ELxZ9nzxpFMzI6+PY+JuUyf82n2w93NnywNIwdWorAgtozbLUT++5Mp9m5kYWA2tNqqi9f4mWJGW
sXCiZmo2cpSooNqSeO1CgqxIMEW1b4VpK0XHusjNhxjcI8JqTXmxkwggQY/Pg6QVMlhK0yiyrMPK
fyxv+N5+M2cl2p95LllHNpf2MjWkGWtPULMlK8E3VWYRXxqLkzhbNfSj/faa8qWtj/hRgSsc8bkF
kdkzkXG3HQSdrJW/3Zl7EgjxgTuIMB4gv5Hdk/RU9XXpZ6/7gH5fK9IyMUzqScWtwb6vUPjU0iqm
+R+Pzwsi+FPi4/H/Y1EWklEhRNfMFSEmDHORvzywCFpoV1JgEaP4KkofIDShUZLz4ZggS7nGHN2O
Wxxk5NrLVfgaotEkt+q5tagaa4OACPWAvuqoTR/6eY2G5iNcxJV84P/67QqkHeAeFMrjDKaxPzdS
YGdNhY5RGDxOGpIR5d2ORquv1rMwU3Lgt3BeXSgI0//r3VmFuY2Wwj2bETxE66eISdcUH6K9KRaa
Fq52G5JuvmNNsrzAIQArrIyiVp5MH1AIyLxLZG6VG38uiCWu7snbRFgY1O0Gvh9WDwIUqSQ5vbw/
cyLOMwWjX59n5/84Q5yvrwAPd1o8Ir2cmNJbqasMJyK93ETti7mjVMDWWMaPM7Et8YNxQWlBwhUQ
qUnblWRwpWCdRJN7HP5j0SNeRgmtfnD6THZN1WPmMaPqT6j3oiM2kRcQy5qkVRKf7rGkY7MK2qsN
JSRUHUQNRjzIi5BycO/DTB1Is1S3mpNX0/gQm0sMYFLn9Hz7qtQC6cVbMPBWn37ViYOd1Mzj/bzm
dR92DwfdR5GRXHBV1mdcgynJ7z8Z575xkcWGCgPdLVD5zzWOCwDgENmEMAI1AHBfMBoMG2lmw0Dp
g6hpgfW52vodHSmxeRReLx8S2RWOQYtcZQtuMMgXkqzuDvJOOl/mgXPnQw0i38kW5wbqxravwNxe
fpcyBhsEzOy8If/k1Z+brUnmYRA7GzZQbw8HpR4hemd4mzp5DBhHjvLi7LFdAngG6vL+cfALW2je
UrBjhByXyXcWaVmbOoBWMq8hb6jPueJEBSC1clPWrYK6LhZDSaxcL/QIxyo0drKYuXKsS+oT8yYJ
GsZYNMZMCj61RzfnEGaRDFjmbHch0LiUhaQ6FQ/9ViCQDpcQPtOG3HfYG3pQVwGehui6aEujCFkl
XUkururHfmNB9LyYmB5s6a6gG4gdnyjY/ReD/QEfArYnVjnxXXJ9S7DnuaZAZ/rXh13nZI3zCtlu
lMfPq1odHlEIy2f/5uWRPcLzc9xvBKYlN04k/jL6GOxFsX4feOxNS5vrEuBkU2sMS/nMGO1zs0AN
PpANbbDWrm+8722BICJZ0UXAdXp/LLyvBL1p5zkhPTjsXgzy/sW8aEco6iTVa4tYRFQnE65BjeeL
STLxsbkgQyKJoGOAnnSg+g+Z7GCVCvwjfgmjNI1q2s7NxJhSGBb9QrQhT59JV1WZReFIpFajsemn
jraqHPcmsaK0uBIvxe7zKhXx8X0EC9UiqPEQZa2TKuNtfbDldfMM5P0pg4UAQSiqEBFL9pLs1nBV
lxePcOGo7jIOA+0Dm0AGFxADsoRSPgfUMRwcl798LkEsaSiRmyKNbuJ6ColdoIPLOtlW6nZTApSt
1uBKMnn1Gn9+SDuXWW9wqGDDSvymyIgH39YkEHjHwAAzWfXsklOMdRDNclNeC+8/2w0o4xx6doLQ
klK52YvnI26SSpx1hX9+1YBEKJ+UXoiYOkNKBdg/Y7VHiQljvm52Oa34tB5gNkzt4wOIjbUyyIwW
xOD2JFq/ESaELw0ebwC9t5iqS7DxBQZTHwYsHxFX7vpJEMtbyBNTBTZOpwq2zM5lODlkFyWm4Saa
1DFx9QNsoJuw/DV0nE8opgjd3E+hW0ufvzgNGHmVTbpYkLaD1lhHlqt7dkxa8WHn7hILxGkpSwUn
ItvvspcafW4jAKvH7XBqWf76xUK/vYV70mbI0ZgJEpon0opQr8GZDGHXKxl2ciOloXaJJgePi2Jo
//KjmdFGlc5LBplpnzrsQGO2UoWZx3RcG8XhfuneKuWZo3DzQBOZeh53ulPfREfjduMgao1x7rJ4
fyOsYnrI5S+htB9Wdw7ZCFR2GYDiFoWvEz5eYGidZQCxp/XfXHG2tBD+TKyKRELsAV2CTd/0u2Un
oUm5EW+v8wgMqi69gUkCv90S7vTA+qlsVu7l8UHQePTEPpvH1LIqial5d5iqknfY/a1zBwUy4xzn
a6o8eZwH0gNBoO6XwVHVnHuX/WS5aWkeMhmqLpYy7K8EIAhkWTfWJwUGpK68u1+A6iQEnpSDcuQm
8DIixuPP8xuh+B7fYWCyiNzp1hmkTyKZu5W3mZqZAnTWVwvkA+F46XzrS/Vlq8C/Fz846iPLjOQi
3PbTCVSeSGj5AQcPl7sUaUHp06ZOC1H7U26idDCcLIpqlH7h86CzoNmfLHR/8C2fP+JdrC6JIx1y
HM6heQsZIT9VA1oRk6hK4y7AoW10UG/KfBkoOPpEWE0w5M6rjhHKGZsxyArc8KxhKVIewSQ9m1yZ
TE6w0Zs1U8Nv/dojQSuZF3kTanHfBJu82JnQCb40Eel8fxLVqDHkLp/AZ2N2s5TTTq2BPkjpvtPH
QgBJsHr9ExwR6y6tHmACFO9iPqxAcwBDuEXFNXOc2vV5XqXmKkpXm/ukfLS5+tRaUZI2ZbcPls1p
0+lt9oT3bf1MSusk+R+0ZXVrJZzupVw1R0khfEwkDBMoFsED30+tgdN9JptmB3aDymwfEh3VP01X
WTo4JidQjFMfYrfImAdOlCyEuq9nF6eoK0F9hM1ka7UeLYaG2kQBWGEuT4LVsMOUZhH0C9hjevQU
88+/QPfaz+mJ+WR/jnmixITDYlO5vfR0kFJaJjf69ukTud0YW1E/CFqJh3ic9EywTqN7AaquKtf0
VoTrii2ZH40rfV80SmGVdIvB+oaefGqvinh8GvzyJOQ7uE3gb1BDCalzJwK5iTcPvBdUUlqtcHtr
+D/x4fmwrf9d4zpqM7vDfQYF1pE+vMXaRrlxqmtLm1X59CuO6HAfoboYVrN1Gp8cUKvAKuK7lHzF
s4N8zKJBgKJg+S6oVZLV2uMcvXGuLPufQICXpeA8laVTUQotlE/XZmThp8civDAk6VzcREUmc7Wo
14vsv12Jtl8x2LUY/kR2igNfOOzDdkBXGs7n2aYPB1kfcvkP1paNN782udHvNWPfjfzaw7ZV4KJp
ylGxi5eDWNIw+a9MDkaopPSz+PYzLXva0WIAMJD5BZXN++KMS3xsNPxGyL575Za1t/B6pQbNyTq4
WqLWElYDpUqNshrTXEc8ATcWKH5Q0ADFvHguo2cTC/ahEjhpjddUhF7OHSlTd6ecUh2BJtwkIzcV
u+1BRrmH+6oSSdBMelnXBTOPEiCQI0AcuWHQj37HwjAv75b88rHgi7Q+IPN2BUE5Ujo7/TRyuG/W
GrJNlsfc0LzEeSHrDcdC3suT6SHsTp4Wa6rpkDa2RhsWFKZy8J5Nw7ENtuNXyc5F6fHAMWdsz6u2
9JDeghFNDj7c2dPlGtkWxVEO1qWfivHV8QAYn0foi4UmlrivvisEVnNtFfaaBKZPPvbLTu04OJpz
/PmZg013UGAi6Z/xQ5HgWNJEhF13vpOQsHgmEQFCGMxBm2l8bDRk9cJKQFfjhtjG/LF3KZcp9nLm
mf2/oKMECUXKW4mI5bJ5vQ9vLevbRwUWhLUIelF7ITWvw5VMhk0Mrz9sj8hhpF7mIlss0up4Uf0w
nwLszzEFuepJaCZi6RLKBQdwnEcwr1qzLDh8MF1Pz/vX0KvkkMU8W6sPFDnRBczNYKhIyx4INWvI
Yk5KIxG3ost9LYutzTsSpSXh2NkBbAqj13jCw9RAu5w9Zrv3UUXuMzHgL5G5sbF687XDIcQDflNu
OIY/xe5ivqATJuL/sRX5cDABf1H+mT8jFnaviyqqER3ceH/nc7y1uwieak/OfgmH/9WOYCSCugIm
P0KSMPh6pmkGtYJRlytQbh6scC4QEdLkBad6ylq46P/QoTA6FmOK9WTij/BylmiNsh0/aZbUoZDz
JB6WRt1Xe63/HDKrQiDzaQDm0n/Lpn0bsXf9TwJ3jW9z8/Tjzeul0cJS5rSh5s6p3C/ZRoRB9UNN
Q8et4WL9bpIuFMNdY7QyUqdCKskPGf3gmealoFeGhWIcpJcRrktphW2TqmygQFg4qYbzAR0FW2Fn
qa84a2oRQw2vm7jJ45e7tOqjuYeNxATFOFZqnFgP+ZQabm47fPeAm1+P6FBdVG/GytuB4gy5bTmH
cqyj1L73L/5KBksMpvBf2pq6DLJZCLS0DELYVJxWjHsbRDnQDU4SEHttA60I/gqxJGHfXFaya1Fo
RyBxYmsSbL2KT4qNpAa4dwVe54frXj1iFSrEXJl5d4xJFTZ4zZtLfPpT+MN+mbneL+0c/NIWEJag
43GOgAX5NQlk69TA2tL/e7jIbn+abG+OIoa9gfVBhzR2EwPVlLjkss3H7+4BxHdh+T6Dw1Vohtwj
XwmIizcNQLQXHtU47c13tS9hSRyevryTBHLYaCpqmasQlbavGA+hAVw0H0fsKk6ju8dYPD8Ed8IA
xKZwdOaYGQJqexWrNUPqL6v1n0DWh5Z9cAe8sRPGM32a1nbvImwM389OwuV6VTKYv/2eq5h7K8Z/
YUc9uSE7mJVyxZA6yH2cRQrAcz1U3joXEy7ZtJyKQeVH1rsOhW6qU8eyCo9+WjLRAlVGR6LWEZ5P
9oeHL/p+SLrvJJJQcmIkuOswR/JjIewK4h4jG+S4W1tlgALaLb0w4/4Z61vRrjfvWoQJHFhACRwi
pLBSxwhVSr568y42qNipvKSqIMvrrrFCP+hMQgJ9D/RuPbY9zg4opQWZjbajMsdVjAB5MJ2leEDJ
0WUJYzJsQ3cEwScop5gx/tP2jLbjEbNbMe3Ka7ChUBVD3NNDwSQ4akfsG12uibxwrTdfBiwIs8q1
4xAvMC3CAqpEsrtdUBeDp+KoM06gz3vcuMJbwUZK3B/5uaZExnM1M2mm3b7u+GIcU0kdfNX+2CY7
74/dj+XC2FnA1QHZjdFkEhBATBNuCwoOsAKGZM8unGd9fiAjumjOvajQNI2kry7ClXdIAcAK91l0
e1mXNL7IGUFJGWcMgM97lW8RB3kPgl7j4MWxahMJtosEzeP3CcC/NeQmXzstcCLEemP7uGqWe/DL
McrA/nueOV5AgNx0uuLrC/Q8ISIeYav57pE2nUU+zhbpYMofNPItz1gVOr4O3zuJ/gFnyz+bcx1h
weKosVrcxo75M5f3RJbAVp66jzpjEupzP8lZqNPNBVP+7qIGQneBonoyV5mRoN9hxzoMjbHgBe0P
Cer87NUBTSWQFJkCv4rmxZzzpUQS6ZEDmko4JO3X1QMr5ngilVFYyiFzY+CG0erfEe3vE1E2PFvf
F7KfXBxMOUVhMh2EL7bk5VO/OvU0SHxEVI6FVIMtO2ChPAJNTWgjFR56NRAScROyduF3iF5A57KA
7gwsWYsxajJQxeyY2iBg7ySming0wU4FFJv6OmeOiG7aQMOggnTxwDY7DONCspt81wXkbz99aMvX
8CRCmGZH7mke1UgoiY8O76MmAblNplhI1e+STD8ptVRl86QzEq18DvXBZZ71BKfTGZ8FqadeofNl
8YAHxbzJ5DiyfWr036yDp3B5rA4hbVpTy5Nt1mlhYwc6Oo1l2TqtVefqGLtIhQ1yGtaz/YV8lO79
zIzLh9EcQDMtfVz2STdwiinZdng2Eq7FLUMyOfba0tkun/w+KmfB8Tnvwz6Fy8TXLe0Eyui9BhDl
vtrfTjoPwCNwt3kB+/trp7nVH43zkWxhhzdZswSZwZU4ONl5tiVDXNa66E/qllSQzO7MlR2sJjEr
qc6rtEghB/jpbiZuUrxpj/rYJNL7GVQrhpEZtDVJSGebmr6FagYjz1TV5lnCF4BSLePDAUWbp4HK
zlFmVwpRiciSJwTjmumMd7ng7KVnpgp25bO9Ifzyw8dgNUBPdU4J1Fgrw2AMcvhKyEjzYpXEBf+c
ydDUf1iLPwFjyWLSJ0kZ65nIyT7qrzIH/GK0rsArggMiva26I4CfJotmRV1WExv2B5g9szA2B/5e
HLyikLvihf2YQYtJ0r9uemkOA74E1e2nM/dVwkz4t47vyPcR4bnTnQhpKCxlIeCMRZstpTjkCfHZ
uI8HpxLjS6M52+2raRMMIM/3kBCiodx9fBv8LNfTBug+mbp62qyP5TpfAVMqImeQBUBgDFK9IguV
JXGtWef2M0q7BHyyAnJlCYj/0GcX97DUAFVv7G35t8E92/FyS9l9y1A2tPsDfv9bEUU2pkjwYV4F
VMjRwyLkIyArDWL3Amlpl40N0aWN9HRPyx1vXlRie8HJ8wzeedYdrBMVKryThqtpYaCUfVRfis3L
sICL5eToBTfNTmQlOKySsWmj5EhblrAE/fegE7Xo64iZYhLhb7uI2Y6oE1H4kNH5xh1OYrwIGEl3
Amtbdas+1NozmXTcq+gajAWNFj0kT/ITnr+sxyTgiCWd793gAEkjWnrJj3twTdW6r+u0g0HQ6Bra
Hzm/b0AwNZwKGjU0yV1J0kC7VkAXccDgSrVcTgrZa+s1HJH0i584UFN112w1jdAUuiPdw1vVgpoG
KVKGLZABFChaXtVw8IK6sU7pi/pg8ZNefcsRr5rcyl2ODai/Wxn4D8eW5Ba6SUTzLSy+o5mmdr/B
27kvlY/kOxjosEOTU2xoJHaBrwNuS+yMYSsqz96YaKyZgtudQt8J5ITgVy9PU+xqzVbgd/jDVtrM
MeGKXxgay/DDT0OEgbk9kVzSohhrzAhd5ArvDGuDj1hpIKDRHPb098YBJaA7uTH07cjfG+gEqTWl
aloWjGYLT2nH/Mdx6QtxI00uwqkuwAYs+M0N2+CQFyhCo+NOJGE8IQH1O2gn6aYF6hYlsZEyhCLq
+YuVMZpm32SqWhwNM4PLsUv7LQlb5QmjS7JT8wJj5BK2fZqYFAGZt6EE4TWMX9ToKQJJ57BbLVG5
l4htEA19fD1xoEQrB/ah3s+3YxggO6b1CJ7eFPgyrGMq5GZt+7mXfZXb9/uF2k0atOTc+GVhr6FU
dniNNb0Rc2me4+y7Hg9pN0C4OZTOkrdKzOi1D2aIOP1olrvtaKRX6Up26wVv3qv2kTYSRQWxfG9B
FHh/iQqZWdNyk8Xr5CTJ+G4UkGIr53gKUQNFBztDT12BZogO0mrvmw+3eHTWzC+uh7i4xKa7AznA
e53tEtGHX6GdLekZXafCJD+nuawGNYyDQhRZavg7EWqQXDEn6A2A/3nog9de/yfeR3ZI4nD+KWuG
enyYyehCVSGaoWZzK/F4CbU98MTIKXkhbUJmJFTrWFpetmaxMHChE/QNynuWfqH+kcCz2glT5x1R
5LAZx1ws2TmeNWh80MkWR6QeZcaiIRJYcJ/i0flzXsxYRVNRPJ0ayZQ9CSK2uR9b2dBEtQ6c+XIz
YqhAmb2/pkH3ITMw9ThP0ruQ07/qsNLKN4iOxSK9iDlUk3Wz+/VAcPGyUWlzMkfDTWDybLVNSYiO
0nvD5GCH/qfoP0rjHjcZ0k8/2HIqMftOjHtQ5aRH02d1O2tqywS5y2LU0QEOeMiyLsOd5pfqtB+6
hQGW+TSrkxZMkks1fotEK8E3C6Pc0jE8LsjzYXuwMzI9FOnuemBeKq7xR058MpfcvPLU1c7K1pw2
6a8JYj4yH6hisKe03AQFg0yqx+dJ4YI3ZmnIZL8VFc4KjrKj3sTJgAyK5J5yU1kOJd1AFxwYl5i4
p2vlydzT5BsdhU8gjFl2Bdf91scZ2UpUFiR4juXKflp91JwRKnS5mcStJiEDov1s7DAw3BZqJIrj
d0dg2YvGa3xFcBHRECQg1UU+CbgUkvobjo7jI1wWLg5ov6SAnAwzwCQAtK7fIVWGVgWF5FM+iJD4
TxislekYs0c35CvGl7+Xt2BHSBebQxz4yOK9J6gTySNr81djqY89A6aTyy6Hug0JWwB6TaOSJBHW
xF0KhkkpDXZHxbES+T8Ezazb1HaW+HKXvquRXmUZ0EH2p30PkV3fnfrhjDwNaTB8Fskoi7O4Pr4I
eCADxIvlvpKEqABhs9yMy1jW1u6L+xviUxlYsUAEZ4U0xgu6X5/a598MJHEf6eqeQq4Su/b9FcC0
nrTKGuF+rcarowM+eA8v7IST2IsN3HRWNTJ6yWDM8CFuhdYGSFtnIUhNmeuzjmwdXRnglZCIXDSc
LHPIN0+BAzejdOijuecmrDc1DWm+iSByX15YUTgf3R7vWf4FSbg7tGfVB7IQM0IJpxiye6EVxSHa
TkEOWSAlL8nggBkQAbYek3AxrI55Tu2CwMRbW3KlwU1i3+Q6L61yKTuXzqGBAkTq9sKtUKiWS3Wp
filRz2zTCA4N0MXzlF3L/bKo56FKRHoi7Ptz8sfGmbBPnUfMUYGLUhFc8/M5R9S0+Jte7CvjIPbL
O/kPoKmZBIEI4Uckgx+tJwwYCvsbqKqayxG8Lq3b/lsZn2jOstTVMlqQi8Oak6x9+MRQSZXN0KQJ
WBUr0V2xhg3U6M4ZmZR5R76AO79GdduihNSECiF7qithGmJ01dOtuwJsdIZIDLm6YI01fEzpgDOa
yYibYTTN+veGFNDStIINSWzMjIoxTV5l8+uT1tnuYNx9FGS/AJtUAgGTvFfGNebdgjNKV9D4IBvc
AbriB+mNTrP5Fif0LIK8nlZCtRaT0MKRCIeIICQurwFbGlj7ousxOaQ02apxnSBunxeFe/dK4TtZ
cr6GHrGALqMTwxGbxImVJkqaS9hDoNCzfw70k2jbpVFJfRfl1uSwWh/iKemdOyOwj27I0tbrT9y9
dhyKSR9q+v0caZPg9kMLDPGZXGZLgla3CJCVjovaIGoxY7IinWAKKcea510CV6fOxGQdwyE9lOg0
vwAw6zDbQJzhuHJbffLYBANbODdy2w+sw0j5uYe9tHWr3z2GF+RP4aIXV0iNHfNknWO68hehTopR
cIv999V6Buqn211Hxz1+BfAHeWXDWJmO6YW0D21CCFtTnflsn91vtaAWsGh8D3hhX/LEDtnyfnlZ
lGBc1/qWfo7X32yZj+TgRnbLwy0r1whW9YntiU1K8Ks8EYmSuqzdW7IgBi0K40wGgwmWH8p3LDLL
0ce9NAWgsNCnpX2KUqQi9vvfZ4Cj5TsgH0PaYcucCX7/AiHWd9vbvL1bOH76N38aVH8giFGzbLx1
5xYxO4b3x6khXGODxYYwyFIUbG2ZQl+8tLIJRQdjFJUCUO+CngU7qz86DmPmOUjaD/G3uIVoUG0x
VmkbO4k/XErPIUeurvdHQwGvpzhXNsNV/lLAa8XMX8QnU/qIeK8LN2mIj2IEuCX4bBdJ9FtKJ2DA
9qy5ZFWfHj4OEwyUt6ly/WexKXESBTX9T5LlBPHSaIegQILrHCm/c1ZCpszUvLDWuCOtqJSn9XHD
KcR+PYqTfyZDtUxiR447baMCPrfLodMfpaq/mkl4v110owwi+l5aAaXQR7QXaQkl52Jw2JwsB+bC
XL/iDAeE0Yn3PHv9mG+hbQCbEe+D0WXmLcc51Dh0E21V5cCoCLQsONeNVLuaNstfZlD5/9NNCsXd
kny4xSzTe52aDPXX06TYIIfwQqgPKc6A/DQVM0/93Cymmh8LTq4nRe/104N6MPBACIEhwu9nPNjV
qXzmRFA3NYCaFUhhO7fOAWynxHKGNdgTjG6aPgWsGoEadGnyc61eKrN/nlk3wldk45bWxmbaXg47
K9HDzlIVYGFzENLSXmOrilnfpnXpoSgtmoh5h/UMjBnh2IA5RQ+ssEDRfIoJ5D1Jbuu8nNN3Nvqh
WTtIZyWZ5oh9U39q/tj8fiVu6TYl0hyxtLE6M7LfvZRPfqKd7/L824JWzYt2MQbr/0chxc3ho0X+
E/o/ewxHUPzBbyVw8vJua3z1aff9FOvDUh+sHk7dkQEzSlqAK9lZKuGWpar8/Ep/78L8792ku/Yk
gNCdL1QxofFbF6qqhl+Et6Ont9mrW61JVxk8cMt/XrUUh1ofZegd9HDkRQ5Z/vx1xzJZiV5S2aK+
iuq2k0/1zFRBML1SjzJsUULPQuiR5G5K8WolaqAV+mtBXqcVqVcQ6N//JnQwjalEi20wX8dzmRqB
IYsM+c9CaNCkNrYr6QCrAyq9M8WVf4tykNu5PbeTdLgmdzuowEMAJVsAjGwcQcuCQzd0Xf+oMuNO
UKcK1/Smxby3zeFOAFeXr54MMUSQWeeJseTbuiYim8amgMOXf8PkljpUAtiL4z6MtEDPSCISmkBc
n3+jYLuo9NnbiJg1s9VDCFbBt/Fuzd07uPm/NDyBa/4Fhy554GR7otWRzsd+bjJIR5qb6+QM7Hux
4cV0IdiN4qqNLaC3w/RF6ryEbQmbbFipwSHANUxDUY54bKZixzlUjMJKG246KvKZi3YL0sJmM/NI
nwNGRAmsr6ew8ZYKKmQnNHFLsTx8vFoDFFgdON4ccxKkFEjSzwLyZAuJO3Zh7HK0HH5VQd5aKMHO
iTAeYZshyeJKRwBphRQK9eBBZxVrlwS2L97x1+bEAfCtldqOiPlqMSbhLirJntB6eynov+6dAm16
k2m9Seegxw/NgLvWxxZled5pJSnrNS48iZx8wC5NcWEkXbY6TU3/83sIEtLlBIBWa/gGvAh84dXE
F8Zlb7JKqKfb2jM82qWXPIk4YYEQFcG3p3gAeHyzIwbaG3D7z9pSfdMXpzJO8GW53jGe3NwEfpwa
UqGCKfsDIQMXYeMjNOsEGgBatU2CE8VFnCe1Ol0DbIsLmKZ2uLFyHY8dfvFk2BEYdHm+FWyE0+mU
F3cdXC2P1dOKZOTo/5HbWOvnfX3uhRBy7OdKuUMW3KWgpbpbu+LxvuA2oSzFXUgu+Dviz2gsEbGD
tzfSVxoXPwDtO4PW0+YMrZ22/qlRIhdPzn+ER1KvgDqoDDQ+NVWqZ2cRtCgNh6jxeTro6W3F37W3
EWSUjCCXa01oF77p4pkzN7Ll16iRI2KEjZ+ezFwO4dJnqi9d9Pt4c2p1EdR/PLZafBroThSU9YFx
q79oRZlGc0sVs5B29e2BARJqEugZTCwF7k/AisDjsTX2WQccYIAzzYjDQehYkPMC8IEL5LqAc7Ha
s+RaDsBK+D8roQm4v7jccrh7khE4bPS7a2Y5eveqixySsYZ4+cqssPbgLJp0fqbFOKbmxGyt+Hf2
MJaFjX4fS498dkwSc+ssNUXS2pFykYzoyvSzj1Fowg1xyctuErijEaBT6rtVghuAzEiObVpqnZYC
eWCDG1QylwT0+FgIi68xhAaLRjJmsT1QUOW5r9csw4+svJs/N8d3sLO30nIdxXNDsF21UGZkSVvG
3WPJKDiyKwZNJ5LV/hoNXbhXzv8OTmvnipy211hueuK8uPccoaK166qPtXv5eD2M1O8ngIwVtKLh
ITQLOSbATQIvrcc9e+Dco5/l2bICMTLY1Ho5W37j4DGXtwJwNCp9EpfJv7tVTc1ktJaP35sjHjoZ
5Sx3op2eY2NzRmmVdR/2B6FqwciZWql2otPJNdAlLCrxeM2npjbZSJnITpH8b4ftnCyfG79uUD0n
dWHGMAYVMX3GMXWAPkZHF5mAABqb9PBZ2TF2BYIJCwbFII+ZVFt0LAN7uKiIPQPeEHKP7LkcnebL
6DJMI5TZmKl9h2VN05YwSbcebrgOsMPtziDYW5eIj+ei10CVHMO+GXxtPz/1y/4q0/NPJPIQztu6
xPloaLzcaZ3ik9tY19YUY7gg7KvlmKOeaHvnYrB08OwebeLzbpzWHi8gha3wXAGg5QGY81Yi7Fso
cyX/dGlzRoZAsA7ybXgGa06UEPc+QowOqKSsZ6PDunXEgSXGSxwh8LEKq0I536yItnE4e7ZwNACb
1KxjZEFVAIhSRULZExG/BQ3Edwn4nmpDUM0ZDSl9UvIuQAGJyBXK+aELzeDtvH/n8NNU8ixzPkeX
daiLLsaTYxAsiVDGflwG4TOubmE4mjphd5PP5QV6vOQD8NK0IiYPyflWjZl1hFhYXmfciXpaWSbV
N3bGxZCA1d/R/cL3AJDVPhuqt1uXm8ZHGWHTKGwnJkWlW7MfmEvNlkYCPAQssmT0YHMq6Z8XQqyj
ULDjDt4o7rO92GYrSWqdOhjyaw6L5rGPrYjso8rZ8wRC6bHjzCURhI1/ovBGMErJUlFFi29RnNEw
I3R7tp5R6/ctHLmLK+4GCk4cSbpM53/RiGo0owIlYVlHZPZvs7o4Asq1XFktPw5H1Ppt9ItqSAsJ
BELeBbvR5Xl/Ko/OIMRlctpRNpPg16Sv4vdaWVntT6jtvjjmCbj4ae08KLRipT5UeF+tCWO/YBNG
BBpKQwTfaQEMvFs+N1s1fx8tDsvrk0Pso4DvU2E/wbcaCtcaq0TJrvim2GWttFlxREhkR7tVnM4n
bb52bWTpn3m/efPTtcJ457/Zmajtgi97Ck0fGxNtcelxsft6ScKPH2XRDoh28mUnAUGuzNFggwfZ
EQ2AGMuDpWSFYTNWmffatBfTbRSi5HkX5Zjl56k407JgdA5IJbdqTGyTyubCfvuzaNJ6hDrMfPUG
K+jequep8d7QyMpXExCMlvpFKin9bYnBldmScOtavOh2NQUKvKNIDk9z5kBJp197fPB5EJYZrq/W
f/AViFQeUtEF3063V8re1ZNKJe113bLCj2aoTXwbFli6jeq86rnMnwmnKq/89BbjCplpI30GapAH
M3mUT9lvfkBvLy7ESJEQsx52s37SiduL1ZUCJGahI9yxklgrtTPnONmN19cfW03Z+WAGb8CgnIOB
1I8bEh9dlDAdv+pB6t0tebSCYOh96EZrazOAVuwv0WYb5TCw9Aa5MWg781J1FP/QsGmqtc5t0Yil
jtmICeLszEq1D0sqlxjhjCQe+VhLjVFeU2skhBPWbXj2ABY9RIQ0vg4D0h5mA1qRAkkYGEB47T6v
0DqpFDMgPE2+GQ5oLOg6R+hrxZAO1um6U3Sm5P7pVSjO8OO/JoLjDO75Ne9HqPtROdqKZAxRHEkI
uAeoomH9msIlM7Kglr9BN+CUkl5CA0QnCP3L18OW/RtsDlkdMrT5XTa49bt0MhUYkGG5eUfSJkPG
TUm4U0of99e8qkF48oXrU85CHlNgLRraq6dfbNNMlE1+fasQZTfYlnP1BfGs7itQNQoqm9M2tp41
hvj5Xpf9hSdLS5itleInju7VqIDLpUn8x5AS7t4gqje0YAK5w6zeqnHhbJmUMBrzF2n3v8eBtqbd
NBJAEYLL/KTa+dETVEsJAloa1fIhssWYJoK6Aofnc84TT97o8pO8+1qAWtk30SW+F63OuxRDaZjg
KlRJEXkFDgmeC64LBHhYVac8TYMKh7QrXboxRZWxBmmGz7p6BZqpFP/JjhguUAlje2CMVZUR/fB8
HvJpRAbx8Do8MVRSAueHPP6OnjtrDjlLFcKWcORtsZXQtSUz5m5JEeP+7SQvXttikhJ7G5tnAsKp
WZI1MaZ1OiqX49DQCzuN2GPI/2YvFvxCyCTcHNk0jbs7lBGgWGOOR3BfOKjm1tB5W+CM0AIXi+23
JbcfUIHu1RlWN1SNtLS72jFYwWOAcUXCxFdkDtjX1Hvb0naCOLcKsWyM/kBJ8Crs/d26HsCJo3kH
LUNjCquStLn4caZi4I8iakyGWwrYiYfDnv0vAtxxDhEp5e9R/XAJpp7dxlgPcXJaO1R4W7jq1Ux5
FZWIDE19P84ldd1uOXxAXecR7ske8l02UaB/R17z5sEg/TUHJmmMB55tncTMGWHwS4MPrzp9aO1J
H5QKZ4ih1eDjIuAG2+/rNiEa1PV26IKvIkDg8fEYk2hOaVm4hMWykGNdZJC/pDzUkOMgmgNG4TmJ
lL7P4nHJb7xqlJiBN4z3VDRGtf9eXIfdvuNhsrBRulY4mhjrJ7hENq869/mtgL4/YjPU1FG06BOO
TpVoqVTZkrluyNerrA09Cy+8FnKGgIHngq3ZdoRdQK1ssnRIFBF+W+snsyBpvx2oLHuww0xoYCDA
jd+F1NFnbl5rNrWAuB2J3LUBTVxPxbbu7Ogosm1cL/qI7QaeTJ2fYL3qg8nVSEtoYvjzCk081M+1
ZnWafWBwHBTABnvczas71lwtUlzCG0QYc3ozEkVN0unb85sCf2qLkHNOp9mRLX6LvVyB1PUxQlzL
X/ouW4Hfn+Af+OmNZofZeQZCBq5Iszc5tB9sc73SZ10PqvM90EltM9hSb09uNP0Uh2HfyLM/d0Ru
hUPHBqWnV0b+MOF3m6Br7gV3JdqkuHNB8cPg7bLb9dWY764u2lOZ5fk0tydibKlN7SgbyosQ9NJB
70Eqh60deLJasHitWeAXyMbqO03F+PKEl5xbaqG9TOnWd+RpuU8HyxIz5MIJjE8lpV+sXD03fkFS
7fspOOCl/DoUVsXBUkZzRyDvgJYMFdV47bAHn5wZbCZ9OXkTw50xl3eHicj7RH7uuQoQXwhAydec
Nr01ihcFiDbeiMdE1om6Fm8r/IdaTAOjcv/JwgobqizRgEMhBsByKPwcoMOIBizwHpV3P8gA8gWc
2kVFOsR0pIFvOXl402MwGTdhVEIvzIMnD0+TAEfKFenZOwnR56glONKqaJkjeHamArHxHT8AYn2j
114paVLqAtE7omtcjjxiIJk50xcEwWcslveiw0DimpquxEDrUdEyTuFo9BDJdHf3OkRNbARooWEB
+Xa3zIXwv2kp+QyY9P06iyzZHVSV/ju6qYPDUzlMYKusjJK5QCUWMaC3GXYzn36LZ2y2a+17wUEX
sl+jpeaPLpl9U9i+2aduH8caAz4/KJXTsXwdIhR0C7EQd9Tp+4b8I9Mzq+jIaZq7KAVOfQCn2XKL
j2UO3wzcXYC9IOevme9VxPbqtMjfdmM41HHgjpMm2xq7cAxVhd5z+nCOhWKvYPJC3m8eO1kqRq8x
N6b/D2F5CT5O3issYdTGTvsHUAlNMXkRuAm3BzMAHObFCF2+hPb8icyMSmuUBwrykLq91lHt/BRP
7dJg+pg7DKH9mlY0rmzk55GTU+CIpBjai55vR7dbGUjctdOwHcH2jVgosmJBa6IlwYcK9kAZowYl
FaGEo/3yHj3LyE4XZGsSmjneL/uXmS8m5ogsmvWDpSELd6i0I/4Gjc3bxo7RPuB6FFQhcIXg2sjx
Mr2cKYn+UK5GpEYdNXS10VsvkUGVQQFbiC2q41TjtYmwIghS9k3en5cQen3Sa2spTKWqWhxwGKu3
nwoEKWGEUEN66IouoNTI4jbtoiUMlRBFhcfpp7ZuGYc2iflw1oyxAyoEtw65jEQ4lMW3bEi/Fi1G
lGllRxcBsqAZmh2SguArUFNehcdta3IDl+hb0ks4xM2m+mFwBnAk3/Qn0SYlpTsA0M/mibF1NIIy
PLKpln+GLSEuTp0xKgrIS/fqb3ApVJOZSO5m0b9TupdwXB9wR57lOSbhYp+zAkWB9JAdPON1h9jM
ZvEbHyudJ2Z2NAW9wKQHpkwPzFvq0UCq67IOabvLMklisg5951a5UHdC3s4+CDwTGOf9cOYlNVMu
tmEtyTAEjfNq2KUUS4RCAmV5gZ4lxjrUmCOHGDpgUHTmYcdLz3527S1o6jzBLYD+Yoaz9TCZxa69
vJBnuIoQsEdirAYKYOX2U2PzRmAhpxWugqHbK1iit0h4PR6P2n0ws8U7OtVAGidzw63DckkTYoHX
5jaK1F7Ky2jaYPwBHaJcC24aCNh8wnxiaviY1LjWZv9NowmjDahqaEEgx2ljHBUE5a5WYfdxuVuU
wNT4brrU+SkfUrDOYA8hY9MnrgV+cbo9CFYZLx0O4EFrMzhkdwAGkpxMYlm+D4kNPJ1T8Dz/1kUc
xh0Do/NFyuKA8vuyI/0bZC7TJAO8EuyHEhr41J2ce97StUUaIXnt9Zva6W6gg5YDBa8hHKoqeTki
CHf6jTQQJNQzPJ8IwmfGOFKUTU8mt7s87/Pecmve+oC/vaqZ7GtkIiKw2HoXfkxPjg8rdwy7HImu
mSNgxCCett5KyEZoEqa3KUpaQcgKLlQLQET4KLiIuodFZNT+mBX6IBsjBCA1NTgIfnaZ4Iu8jKhG
ij5SMl/4NCaWlitkf15KNtsroLyw07mZxVFQ9SgMsdCV1aaysI47ofkLM0gHRRL+Qp0e9xslGa5p
23LyIyac7TjkOInoR+6vLG6P39BPUkfstdTqiS07denhfPwksNl/Bj1lq/jB5r4jqr06bPvDBNw0
Or5hCPD1/xsNDAYEEpHrtOqCxU7sYdccgWqZ1vj91yJez7yCfcZ3e8CaNXircgXtiKG9FW6dWtsw
z3x/wmhpne8hEKqbGvSAT056RVDh3Xw5JeCkBR83GMlCrRTwDDFioo0vskzv61bu7K/E0Pv6pBKG
Ln1al06Awwk8MMHe9W/WDCnWPLeW0E9COC0IhWDe6u+P9F3qgsaLWFoGd9lF1zPd1s1M9hm3ToqM
g0aUmdly0AP5gqksVEVr0joOks0dgdPO9Ev4qesemEGu/U9RL9qHR95VGeD74Reir99KFc/bKiRX
rNh7ic+nAJPw7If5jbsW5WjMlWLjTzEm8iMNXsuUjCCY9WiewpXQwd7OQYnJy+CkdbyJcoIPiJPR
z3u9J6dqA7uj+hchb0f9MmLEbq+HIY/zo/bo8SphDki1Ul+XHJFNRGUnmaxGCL8090VjbozBHVCT
c7K1s8vj6PH3pyADJDeM8Df6ael34hpc4OBF6oMRBN+mS1cQCzKHDrM3L04/bLQY16f8VCYPMM/+
XZx6phzzUvkq6BFyAz6OH75oNNm2q7cCa13WdbaQoes9txfZCx/yWnwYB6OZCPUOtjH15PXQJclk
nqd54yRIn9ABEPr3sLNA8/FQgsqPTG8ZlMZypSAk9+dZ4TLy2CVKm5kc9KUvkE9r7gQWV2F31L0s
EhnSAVrVsmYQCJglavKbVziJqN9L6BG9dAtObkM1cAC+xVXkVW6uLAR2sAxVMUaLv8BN+rJ+9khq
L88771olgYJsqVDuREPpFTIwMbLrwgBnew546khDlIpPrIkfxbxKrIGTJqwgdiiOWw0GRZe8ojSS
rswneuFjloJnOq3IyZp3Yv8tUPjXx5UE7HrEbzqWiqckGGv9/a0+oA6SP2APQsjGsW6r3hyROjsr
hpule7X0XKrrYbJh5qO1H3YYaA1VVNjq2RNYcIvwNqEbTAjPuXWO6F8Q4+QMO4ltLtR7UrO2tB54
N+igdDMJgwhkJN3hKc/k+Snt9j4lzxGjsaPq/nYWkCPmay8yct9jmfQ9rsPiAelzHls+Jx13Ux2D
Z3vcwISJVwRvR/T4eDne4AMT3AFqMZMbQeTK5FYDxg5fHRcvQNxaPV/AY+2HPmNdbVw1FBr8JYdG
iWDmmgZvmhTVjPKOm4n2jFRL8oGg5ashPBZrMp7ttWvJZrOGdgKWKbGxTxpC42wCEiI8UQcB7qVk
dgICljMIAXlc506/izcAKBy1aU/ebR6raI8zF8UJPvUA3WcEMZAa4Gffjr5Dbe+TyR32ZmTddJx6
wV/LLPAHXEN32LYTTo5hbVfAwXj6ic7+aUebYI4j64untV7Ka7Jyor0ck+Fm5viOsDl5M5hOv17M
azbv+BIwQPWI08jx7OUP62ufR0RFpqudxKOm9YcYVHyfeeNFf0uwuXAzhdNDNcZ4ShOgAPT5QWpU
S9s6Hu0+rM0vkscyVrYv9ay46NFosCC+InBpLLfZ0U5lEMZjQdBCJlxi5CUMNUWRZmtJj7kcoxQk
XlM+2VseIx9+D+l591F/I63BSYDdXae4QP7QXbiMkVZz79czVx47Czp/G69ia47TvSgHf6mmXfnb
yEN+JV63fxXDYmH6D37AavL/RXw20bKsngijxVcuDCA3GVUKOqOzYP+Mb1XGPFBTftUzY+98yCKe
CiSvq4IjDYZiK3/FMp3n0oZo4q3xTVSVdmI6JTTHUpWJtbtIq3Mfp33/7iYjIaLWJE6CghbIfx2k
BvZ1QSeQ9Mu3soV94oLRkUTb18w81HbPjEPIzWdwMqhTRYUehpjfaXGrSRw/KG9o6u/0teYAAOId
PGKaccCM5j/M97oWr+eCnon0Q7MiLojafPEU+m//q8VR12jZahhTkaFMl3KzUARbWc7EpBabT6Vm
4wK5zaPrXpG1PQabKdEMc3ugOsSr/V4TWjwEBYgJR0Vwkkh2PcPW1S9g2ceaA2MQPnX9w/5+AHf4
gErPHOeGLLD5mgHNeV1ngMxX3kESgNu1Y8lrsxX8ButnbWp+IaM487vF1ZlSDEVkimWYGCZkKZYo
JEodn5ul5Hs6QJ0uARtrYvUIaHROv77yTq9AX2eWRp5VNFPRlUPGZmo0CE/TrRZfZoaqRytt50NN
cY3ZctCydHT+im/uVHEA++ySN3lTlgbOsp74AkE3uahbkohqZBgH+VVfqYV2zASjTy1tGwGMDq4W
auC+MFLjx+FxU2MkRQ/MqvWHP/bijtnKmMG7EEww+rlWCscFc5/blt2sJuXhUIAT9cXLCvLtDboI
+huaOKaPBT1Vp8dLvGgxNZ2BLxil3EGXsqyYduEISPpN3JrdwWUZC46AuCfA5mVtnUxSUcpHyCxR
qFIAYg4BBUdCz1SpKBxrK2H/KZpRmDU14o9iHVjkehv2XE93I2Tio7HiqCMYAnehgOYbnHHb5Qz6
K8XzHp67cp6BDOtUDt6srHyc2JWwp5fgj0PORFHkVk3duglUbh9Bb3Dg6WNpvXnYBX6RpxOmm5zI
I3lavaewOg4ELO/Huhpt0xO59ZaBGyL5/Cagi5Q1LbQsfEB4eX4Di3Wmc9NsHIW7qAshHdF1tFsQ
x/5nzNrsZurwsVaWvz3E2Car4n9BVX4vJD5ujA5DLkoKuP8aqJJxPa4dBP0TPKlQAZJO2Dou/qlb
fNPhHjrTkslJKgisU62UOq0QSO9DSY3rn8WAzC3bbvFJtRGc7Jbu8lustY5GOAeMRZH0yWNFjHW+
u1wAwX3e72/RzYmcDBNyXFdRcwXlz3zpBqnTGFr2kudag+NUBfm5MCap1DiOJLnNMnrc6sOb9Bvq
vMNZDGBP1vdBoBG2S0Hpr5aRbIRHG69639kN2VPd0Z8IToKdNTWR5eaSruoh1CA2YC5bSDE8idpg
2gX5mIn+oSGPBt5qBoe1nHXtDvXltQ8uq7guI5qDCmRFo2pPW8x0L50t7FNnBRljJpboA8xZGpbo
0Gz0N+14RiCpOn5SlnoRMG+7LFnxjLnIB0C+svWtakpuOOf7gun69VoZ+WakmujeyPQgL8Gk/mty
TfWJ1hIPsd26e7NWj787/OxpW6gGiEFm0/MNF7Qps7B5iULqeBbUtEB0kbTVEFD9vOiLiaAdQUzs
yPXO68PiXnaqIV6wrwSX6zJ+pWjcO4Tku0sSHIfaOAP0F/PAWH4IS4gGgXL6JFxcVra8GEFA0GIl
z4NLMGKxrn0nXvJxD5vyXHUsbDT6hpK2rcUwJwd/z9ChyUPgYD22dMgkAHCqTX79H46fasypDW1U
G7km+LRY/NDgOWDp0VglZ1o6LyU+Hrvya6f4J8k/eNuk4SbgDx1QDIib88tpVNvrvQHXJ2xwUfcv
gIc2ZbzIQ1M831kur1BRUp92BCZ+mdgRSx+uGQ5IAGLPvFxFn5Qckr1d/F27d998926X4dcWt5vV
jtIkqxUuJRxOsrqt6Iatng7tdPfvyALKSx0ciFbYmWlh/BN/8DeAwTGUYQMnyXeteEDZTKAwEOOq
DEQRuhrhC58fYyHTElJK0MfOA7Qh3PBVBMaKRffdwEgYAqQefwxupxf77/KHOUzcTDL0IlKtRlgp
RTKU5hbaLa1yoae36vwIN9BN1veSxAuRU13Km+besPpS0IK4GXE5T2QN8UykoTYSmc4uuOmbMx0L
7BQYtuOWHOQeAGsOUmDD7oXbCkSW8BDStX9gazlOg2UiWdMrqn3gZ4T2YycRF5mrYG2kcSGJRlKL
TPI1p8CsBT/L81/2vMdNoYMKNjz2ewCT5G9MdS49khIl1S3KHp1IvAc12YlqjvidAo/+5fhF1stm
kWd5vRF4fgE3eyhY04zvTiXI3UWVG3gpi+9CXmptzjNhUsx2Rvjgc+iCu3CskuLoDBCwj9hwARX8
LaX7OihoBTo22d5Wo5Y4MQalgzoEtypL4TLQUZ1R4jNOfviUSNhiZdhduR7qXsahJ1Q6iU7OfC6o
0PcxF2LUkUurGNjU6nFeDi+VHmS79hW1E4lkHA49DJmEOvec0WxBza4taluRjL2cb7M7WQ1+8FJH
p0meetjuCODURvwVRgdUCzkb/QddgXsBVBhWguxbxumr1qkYsZG/UY7ipbiICNiDLpiRONr3zCJW
J2Xi0MqE0hJteFU5l+Cp3l/wTU4XuNYlJiA7y+gL4xXugcZs2nPjZLRFVUxTsmy1liByum0iAX95
VHRPuTCsxklZhuFH1jfVQ2lV+rzOPlcOs/VMSFApCqc+lZuzMqvSjOvZgsEP6TwfdzTvhRWArHao
4Xhv7GXId+Sefgf7Y6dLb3KhMfj7LyqblHclqjEgNZ4ahkLGr59xAANsZTyEESYLuom9VPVAEIkK
3U5e9QQzNQjv6PTEnwd4Y+H2okl5Z1pV5gncAuO7H8CFaT2iofItGVk7u5Px47IIMI/els8aXfrE
QC8+cQ63sooE7IQ540WgHoS5IPyEjSOuE4Sp1H5pMLF4GFHBloWr+2vVL9AqMNGpkzXJtLDuEhqL
xZfO3YHwCnxt9ZKC70gO39XPtZJtzRcEmzB+1gLMjYG4i5U86RWnsOQlAjG7hnEIWlvTgEwAotTj
/IhFVcxAj+2X7G//5xF2fRq6Y9CiNhhzKZI+Cn/opTM5N+5usfjIetBE2cJPf1MBHOhqq4g2om7U
QnHDytZsHiZrQgW1hQHrUhijDBsQoPqkyeMyt6nvb1bkjyOiCRsH7cKx7I5gVRkh+o7PZRjrC5/5
cJpYxpzA43nAGdWMJJ2niu+DqG70aiQGTX6vt+CykYNo9Rw08rnZNVYYTA4dK6c08TSiQ0Vxad0X
gjVSTCgwki6Mgcq04gUUrsMh8ODVQpMPlgGb7f/8ywYPBeXKSXz3CFRqgqxrBJWPTEio6k1KVtwX
OfRha+Kl7ZV6YC1L/tnKxSbxnOVdF9JWR8Ued1CoP0tqD/m50g+S0gQubOzB+p73LAp4dKU32Dym
xKzf7h3PQ7qu4sVlHzttfrR/nxV/YBkDF0sjp4yv/Z5or3dDlTSz1tTxLkd0bcUM7rG+vnLLVbSn
DRu2eyWLzegFyL2lkKFeQp/FeYzTF7mBodHY4nzO3tVSkHLvSmwtdxr8xldi81mLWeKpIXNVPP6T
DRTMKkCC/qVLVhL+vABq4kj1jqPIESRTKDsodM30XsFdwwki7TxRfMM8q2ZsO82skZaHGrUNilrL
n17VI7qCsDrIaLlE5PVA6UdY2BJA//ZDJzg3+ImDCIR7LoFvGSoyRKhqyaqRjCeptqKUY5jAHP3p
ZiMkQ9+4m9zubIGAeH74Da0V+gzG/kmlmUeMU4YczF4gwYBuGOmrZitPsnV3s2FI0VHp0vWKtsEQ
zdxmHtKwi2nSwCBH/iXMjfLruFFZFEGNUIb+dgzu6WcQiEMKm/dLRD6g5wpXai7iHRsmNJPsjW2g
nyAOavxF/Xn63/MTUFva3bb3pMG+lDHFFQHm0eMEs9zxc67eP0i4AbU/fKQ7m/YKnzBu6QwpKxP5
wkGzCv1pzf+NVnwoZFUb2ausWQGNKtwVFHbkBqsfi2Pzfy0eLTtFrlRfo9Ao4c6Js0CnXMcCROMV
cor4wljJ5ak5/WM4VKz1IDpUz+PmRX3OA9Q4WjUanjzIj6aYc566Sw5FQpWmexJHh8NsOTW9DHcS
LltCRVfX8WfISuEHOYFa35TKTZRGzdho4sbeYhFCWc2nqY2Kd/ceBmRXnjdEnl3a1EReFgd1aAzh
iKQ4edotp2y7rj6/nXiHlXWobLcDOxHOVMd1341JhG4rKJu6yveWFzdVjXp7M9vocrR++zKV51s/
Nza1+JjRknV7bdSiBCaDFUY0NE99p9QFfvp4I47/zhiXwxksr297wNcwKJaDVkIzs6YFkPzQraA7
iHdSKdQq2hTea8buub6GKlcukcxFX2aQRC7udA5btwFqtk3lMY24zuFpS9qOWABJtFZwmb8xw6Ev
8f+SFnY5Sc5lQaQmCjaj6LsVBhiLNTmMKpQ32gd4HAlkpZ0+SZEjSh4qapEBL3c35a3N7rCXv68O
8GWei03tqXoaMRrZQ4oI45dvkIGcpeT5aNZfz9sw3MsLG69nFGjq6MVvfpfwJijPIKcI8Ez3dzwC
rKw5VIpE75u3aLv18eYjHkuwZkBSAGUHUnkG4xIFyHJZxeEP4fs8icnMxEgRT216XD2HLgxca2Tg
AykNBCwODQlj7jcY39A9TNvsHMp/AT4b9Xg1Vl7UVNDdcOjf4A0C+Lq62aAxjmRDTKtY6q7HTjmo
blnVFg2fpOjz5VuW3JzEdzrScDvNqW50hLy4vBxnjeNgOL7ljvZIDl7VLRMG420ZnMCONsZ7Us+i
+40lKl+JSwiYr8ihleyj/BK6sW0yzp2Jv9zcb6+OgIOrY8VgXRJj4nCCHwV/soqzqjG0gvisQV9i
dwiv84GdwbnfwYB0e4cAGElmJn78Hqkv7mmms/TPNBkOKZi+dFjVYs7jBHN7+6h6gbhHfidvR9jE
wQfWMzGukaVvZDgHyNylqVHfXkZyCrGdqkTYmdxxAS0V7gWCSwWDEYYwjNJFzLdGv1BeynYGaj/B
yK/Cl5/GS1YpkHDe6hl47yUlP4fqqTsHDok/Owouj/a9OPEmWVY78O1GH/FCsyn46JWIG210xqqe
Zxqw3Z9/mzzGhxjAqV8cYkhxbts1rSf1ccbSv9E34frxSp7V//kkmStl99IaIDK11Gh7lSQwwkJl
pkcDY3pLUDNNvUJW6U/j66L11wvTWgOB3I4FJ9v+Ar1lDsoQvZXLVyC+Hm4OC5HaG8zpoKVsjP1Z
nPcrBhiai2fqUGxdzi+INWGmoVqnpggVVSmW+G8V8bWOfJ70bQSAE2KO5O3WF7zLYZZq4BPlatjU
StLS3qwJCbMFIdgFtYhr0gWlLpdSPYBWrVpxKu3lNb+5aPUp6XMA5yvXdbzErRcWdvLyIUL2vB+e
16P6HaIUcLWrYcqFLd3IF01Ffv5CToiqSZgEjqmVzlZF0SGQYPFgXuQ6dGfUddwPWr6rdO1qDYet
2dq8L+Zd9InNqYXeTrwqCD6m2/wGUZ6YR/yfow2ifPAnZS5dsXVfINMLAdmeqTYnctK2ALhM43nJ
3x8QMGQW1hYnCqb4zLoQTZF1Uysp/es2Q3FIafepsO6faf/I601LN27uiyzyRfsMRo4sXpgfbEjk
KfknjB7fgWNyzKeuA0nERalAsRkQtzWBIEKVV+hLQf+OGhDb3YvR1czw9Kb4TDxkGgXpK+Hs2Gw7
76Vz6kGqqbC1ViY90VSSe1sN/vFJdG3nN9LO/5YErsG9Xc9r5yLfKoDc/z80t5tRzVHV79baZKmV
KcMpL981r+eTkA9YdP1J9rBLkr4xTWAUvH4ngSEA69TQIZIlvmjynxArhXqd8UAnXE3hiV02rLyr
hNjBYBhw8K2cL/eoGmJxlBsC5CrlKxYaqzhEnYAKnMDS2u4GUDdjxM+eBsZE0TF4b2HAbct6g7Bg
Iz7Pwhl1L00aH2yVj2CDprCnILUWFxiMi+1v0A2+6tse4S9hN7OepJf50O9yvPOAz/sCJ7QXgB1b
5hBtJExZpYz8hxTqIKrduMyLqZP4wtEzEePOTzSc6776E2S94EoSKCgs9OyIYj8VhgmWYcfm55cI
R/lVgQX9St/1nLLGD/627uvj6AaV6tXSRplJUSkrLBPElJaGWRRUluJlZAK2vBIOkQ3VaDAMbLg/
eE2cxIoRtYzo/pxD8O2O6Ph2YeHURAZkfNL7vrXumJcaAfkUP5lA46RL1twaAt1r4/ER7rCwkxFe
txI1+iWBTAj4k2Wktw0KcKuaXY6XsYY1MLe4VfOD1m5r4nRp5ODy9OID2EYLM84CTUYlUoDnLEAt
cuM8B9EIt0bWt7FwwQXdfCc2BcjwY5w0M0XzMOoOF/tTsMo301XuVgGlrbHp3+k6OOkdY2I+7YQd
rWMG/4AZdnNYpGUhVhGe0PuHb/Y01Vn1yH9gRJJKXxxdiPD7ZjRCR/JkQqLmT9t1wbcbjv/u1Jm5
7WZ3MGi5SgW1ki+JGXlKhkrlKA1OQWGOP2mdM5I0SzkcITwzbXhNuLLq9Eqs1loL72Gk+/Z1z/jA
nAsgQPmqJhuWuAwamR6gsFE6t+FXH/5eSr9ud1X9y9v2GENS80q0i89Wfu3k7sYZgYN7JpuA9FlS
iI/+LT1/jL4IM/MWNXP9JuiChnb7IRJKxKnM23hD/t6S6jgbrvl98JdN17MKPYURRAzj+FY0RUbU
HgTVOVwjXFwMw7ORwbamv+noEXLQL/MJCax7MvgtmyHE9trdi3GD4kYPy26YiGl1ju9yXPksUi+5
Evm8z32Rqrfkm+1JaTh/0ubZlZL35RMP2jktE/TA4zgxev7pYCHzKNokukrwR1d+XTQw0bnj71oG
V+KvfaSCwjCBV7Szld3vi6V+Xk2sJHuoGNRygW+ri5b0BD+cdgUk+UTbblyF/nThkZW3xKriuwb2
LsPFo1xgLpncjq3MbPYJm3RS02S/1Zd0Lbxlcw+965yUYAS4Hc9zHE5ZuBIVal6Dcvy0h5+6FPIk
An85I+7gYknlZM5MCd/jMmk8o4lBWoMi7lK79MYRP8eTIc+YCSZe5OhPvntUcX8c4dPMSRX9zxfd
quKg2Sl2HawL1Oqwu1AzNSQ+UKg0w/80n0JY+RUM/2lH7rkqYQW7CESYZ6HqmshYl2FjgLmpt0FA
6skXaFwzU9jm35Msq0luBm8J5QLl3EUN/Sqe9zBLuUs++UkG2T97ceBwZrjgqQnG3hkkodGW8ek6
AZs+PxGH9LFdFfW3n9pyoPErdDF6HOKQ0eIoT2jUAr7rGDbaLBSLkbK2Qt6X/XfilwnzVv4S/+rT
VXAA14TdY9pN8mBAA/AY8s20wVtFby5dXvmHX3VqYsB1CBPkMWpThjEfL0Cv3VlW0fkDQR6UTPwx
Msm5TtA95BH/57dMIA/CDr9yigHGcsbD2vl4A4CScNuovmc8licOqmkxzbcBDiHToypz3JpfzXbo
gxZLvkqvdNAQj/QX9dAJZkeZ4AMykfFVaJq4KdXaZatU8a2Iq+TwQJY4SZWnkO6Z6h61q/M7QGWk
HRGJK5BKSbMDwtW2WS6U1WaRUm2cgyLMzBBZuIj/iap7IwXFkJXpVqhD+g29Zplh/M/QvjXb77/r
3Zoa18Ez5LejdNh50uOfwcKM9goOLjczhD2iijfji/1XObzcnS/VoDGie+JOKjuW5d1ZcV08P/uh
7ADFUBjx0yqre6uMCtgFk/Tp0asLIYyr349dS/N1lQqOVeAFUisbjxfKKyi9W+ZnXNc6QahXr2+W
VZmpcvpY8jxKacfdO99Gg+P1DrOvDDOp+UAciO1U6L2a+3d5f0m5a6ItZqVHki8rGqL11isBVODv
UrZGm0lzInOVVbusDHCQEwmNywfxN7ThNtupoof0Ti0vaVo+rEF7zJZ+/JxEvhOqSpQfp4EMeOZi
pCkHKentF1QleICMq/5UXYkGyoSdH1iT6Lz+aur+GWP4P1sL+/IPZ0H19fv3KygMwDEQ+SkpzaZh
GlGLak7fvxVVCUHxTvZEPgxYAVTvR3GWVhzVV7AlVQa1CYFOcYoEq7ii0K5nw4IcDAmuMa8jEklm
WaHC+9I4NYSpvTD0Zl4lwpSYRQ1N/ut/Pyha1iLZkX/yRrg6HWwP7ubXGciZwCfAyDGboJ3JrM2e
o35OeX4rHf/2nci5rJqfMdkf7uLLli+oikaOUvnF+xljoIu3pWyZRiCbLAQlgY/SE/M/rZuqaPOd
9bVaL3cB70hYRA/0yUxPmgCLBzTw0do3A56WoKeFLYa5dNHM/p1VHEfY9Qnt3pGyo/zosty3q4GQ
AEuXIs2JUt4CQmz0If4JoLSgFUUUnBhiwQLWVUYieNN6dL6i1kA0grJ/GY7SnDhvH3snIz30r3b3
FwFFpTp7Tf/kLFmsjhIlJo/dk9y0oxd3Llzf76vleIWiSgMAtVbtoD2SRlRlMguYs8XO1Krl+VDZ
bRGA0GzuIoJ68oZ0dNwxwZcXYXItpCZ5000BvLm4G11McAaNbKkadE12MinluUNzDmhaGNX7bNel
+H7ghyxN5yOrUhPHy8wYmBXwSUfU1hfSYqe08s6w2I3pHZjVLcpQsKx0dN/otuud3HtrztbGOO9T
YKn0eLsLxpKRrBnQzu+zBHkr7SjoH7RhqNsBshvZ6WwH6/elQwvOarxxKitKpgYEFPHXfaqAcR/W
R3HMHelc8AmnAHGBt6HznCRVlb9TuXYV2nI7wotKSGWhXy/dy7sILWxGHbtGGUlUyHOdv9oX2dzh
DdDST+90N7UAbL5OGKrIPo4zFw+E4OefaYeltTGZmVJb+dZic5Ohulj3YbWnO06csk6pleE4rnTj
pyUnB1QvrVCakgzNgyxeC9IDW1l5ffIfl0tsjv4Eul+PMAOxTU8nPbQezsoljJ6MeafvXNXAdxK0
yoJCulQ6DUqHdcIYSGkMqWRD/HtybAUrteML5xOpusCsEOP8ps4AqbhW/8gbx2OW13dxTpYwKk+e
NcXdO8MVM3rrH+iN05mgWpv2j0pSW1hA58haE41oLQ3/bbFX1ccFBEQLaUylPE34pdn6acFEWmx5
UcEPe81k2Nz75w+84q/5KS5cIT0Cb1xigMl4/wINLkn3+zIkGY+luWri/gfQvokPIgPFjaeKd53I
i6hY1EPwnPe1XS+01QVsQVeTulDAq+nKUM3vmlGMmg+0MeFg473J+Kj/hWCpQ8+jJO3ClFzmj5ph
xuZR21K0ERX/0EaZcU5kziaZRfj1eEYAENgbbuwy8jpDMEPLHCZBpBAfXEuupPcnX2oBXifRkUrg
aEoRPnqI8F3+9y3XkzNNr25MoB8fdd/LdEgVaUBEF6QF5fspC7okiVnYLaOu7jUJ31lRr9sFvS4R
NyaF15fb64xK8HlWitrY5NLQh/Ihq2oiLjNEuVUAw5HWkdZiwLj91C5oh3DmNnHMPjv2sOvWrgfE
mRFEcB2/W2ybxQV3dS4nUH6/I/cJ9t1+MWD8o+QpHMgFOs3XUq/lv+wplkzlHbn0/3cFioYc6KtT
XqAn2xXjQNmjhvVwxGx31e/l3HnKUY2iee53bEYufQaCk3BN8DmRy/996YxX/VTlKYMWpze+uGyh
A2DOJ3tFXZOQr8MrJS0W5IwAVA91sEBL6yOybHiHieFcG7/CB96/mO/xneJSg8QTSz5CqE7Z/z4S
RchN0Xs0sOO7t4IBgFeyo3QbDwuF169+sLFwXGtFBzppvH8j5eDxPM3qg5tDbvyV2pDtxiDaGNlV
jdPPydbywiZ46BDTrGo58qIiHP8/yghD6sPQM12MUbg1uwMvv/qC0B8o6FzFIZ/kr1eeI39JmjMd
kHWFlnkkp3LZ2/H2JHQHpzYUyCoNYHBxTnpWnYirmVXzXV6yrp3dT5mnoWaF2pqUr+yTk+gxlpsD
neVfzHc4b1JWPNlQDK2o7kaC9vwGNRlQf0YlrIV0ORQTCVH8P3gNKiOXPZwifR0TrVVJabe1mBui
Sj/1v8C/DfUCNwxRsP/DxUZ6jCEFvpVEiEmThKUyNxFJKSw+jYjFwmzQ8wg/t20vhGz7FpcQjuS1
HC600DYoI5CBGIjUycG7fa/0dCnCdsga4+FySKh6gC7GSNTX/rzCFGAAbc0/ywdu1UNv+v1BSku8
yj/FcLUL1vQIIVhfPKT2Cmf1yxyPdWtV4PE30dlah3r1+Gn88M4UHOatGu+UoqfL90zkbFJ0srAf
edTimjeTk8ljNx9uHy1cnQBnid78mb6ca2RnKTC30YRzRpfp3pfvMTMdMV3MGA+0qJYaV7T7gRbY
dAKo5GLzzq2LXFROW/zekDn8/ThYHkJKyQeQoNW1febqy9myQRWrbaalBh22bpDrapU/NO7FjpyR
wDxFnMA6wFtTZ4W1ImCETVFeQPXnSO+JSVyt6B3SvClLcYw8JJ7CaVkFWN0VGgSxhZjmMiJGDQT6
OkNKrGcY6/GcgLtn5OoeHJ25z+/Csxi5BUgEa/0+iP6dboQ1+m/gfV2LUTtEJNg4pDIob73CSVyY
sGPTHTnV1tZCln1S3TXGZDxvsNpH9s28dncHrLAgAnjtofOO+R0qTKRLQDWRkW6Yo2/I6WQmT2bW
SfptB6NnkwFMb9wRpb/8MPe5Ia/fMBN/nPOTfz3L71241YSC2xJwxp9a3M1PzjxFH959tTpdcYav
wDO/KVBYS7qHFRc7OBwNRv1N8/2AyTZGYumB9JX+XNHOP5uaMX4aYFMUHJCW1CKpR9bO9V7lEwUI
8tEYTnVn6XJVqlHMiqBrn/9MUZKzUNhOq99Q02rDhORV+5hRmSWgqfexszXGRjmd0+jhcHmpuqiB
og8NiU77mzAGfenc5ncMVTxoUzRrsBqIQk4dbgwJ7IxUe9QVzt7/Jt9kLNvb4RXmddrKlAtJvOd4
kzwMKGbGvhhNDd1y70MzOGBwI++9E2E3AXw0PA6pxh8KMxQ0w+KpD5NBh1DugQGBdLcLKq0YzP8u
DiYZk6dtisWr63dzUItmuuo6rAsgf2xqg1+g1P36ZAl8PqrsAuugvbDCK2B3NwAoyJc46npSWFyx
pjRX5oexwEtrCiSSNu6vcZVMx3LKFqu0UswELLy61rgoe/tEl+hCsTrMj9sVpJMpzEwDWll4w+Xd
9FokdQPmKdJBHBjC0uSBIUqyXybWZ7k4IbYIXZOmIWXyPWq97/l+PjULPsJRJi+E29lKRqC77ZOI
1dquRlzZffAO525qUXRdCq2i/BZ5TdbdI/wTqVOyFikztQGqGVQP0m9TOf6CPxCChEokMTO35V70
CbjmPY2AvSXRMyMSw/KdxgBFeRLDiLaCrVMi6wVAaDqIJw/KfFWVqnZIOAHC0EXQsEHOuij1ftLH
tUwzbyJc4wG4e+G5dhrN975jEnewHmMNPYdgZ0Sw8xOe+4Th2zStZ63WJ002+zb5RKfE/G3zpgBy
GF5LdT5nJ8RLkgh95J7vjE1/A/H1gMB3fNAsfDmvojFyialg1n6v8Z9Yx6G6F3Y3vsoSKO3/ccBf
8XE7krgd0djZMW1LKl7DN1JCu1JqEBJdZe4cTsBqlQ74PSQwJhInhTSL1HmiwPXp/XKMbZAFYLbu
nVkordDnr7Dj3vKNkuSd/lc7y7bfkT4o8KuueBQvOsUXQTGk5sRESW01o5Ip5ix+B4QlLZiVF9zF
EBrcQ95e+OIjgA90zPcs5V9cbZhHm6srC13ONqFeqJ3GnCzNQHg6EaeL9xXuVhk2qnr7uaz/uO5f
SqnFdADDjLXJJfWzW7gh4RG5TVcOjq/WHwcQWQdlKy6fSECy0QlnN6zIAsx0oQkvQOz+3uUcSnRB
AspLRTecWZ5rysjgIlpHTGExRjKAclcoqY+p+dp56yN4T2Z9fe4iN76QLqNzrctU72aUVvcNmyIN
5xvRWXOA8HRm+wT3QIX6aL/TUdvnXjZmyj3pfhjkDCX1H3uqbuEG5Dxx9uom+7cLvZXxGHgxF8Fq
b7q/q8MM0lvWr5AUIeWSvmXm57LqRcCAZ9PfPrhW2ON4wvzIPdEn4boXxW85YOjFYeh8rTEk/HPB
MT6CmAg8DOOBkosX+MOhkw+vWFrdZHPu+fKo/WksUkz8kVdR9NR6AVAFe5zdfN1XkWstT7Y439V/
xCKdxbFzm1otm/IDJhItLqGnS9GMZtIjclFBO5kzCnHgC6bbRMGMNX7eQALYAHJlbi+dsZL18TOv
6SSzSPfeRMgrFNPVkQplKqkGAUGAfoUT3S0E9aPKHhYQdSCkmDiGg7avQ4DduUV/Ki5FQyujGI3b
1jWkpfkyaZ0T7y1cL6029+/j0EewgW8BYGwKFuOPECpwm20W66M4jFQXbiPcFMgtAU24qlroxs0V
hIwP2g3r68ylwy2J5DulOxrVMYCEbotVEEBvr+wdbAQQCpULujxS2vlfuOR0LZp8sPsyfuYi+0d6
u+2qeagAEe7X8xFvVvlyqZJhhsWBLA1Mvc7VBxVHTFS4pkF966TMV6UL2WH1dzggtw9gZZHK7tGP
itD1PN9mv6LEmRJT0JNbBzGaTuGZ1JNBcfMvLTCzhfHrXCEXjNHMaHHmwOkaJmY6aLXsRdSKW91e
o+aGrQdttTOEWQwmy7M/jof1piUfg9ezkFcuV/rdv84/TyTetUdjSIofvZ8VHIKbel7pYY9KV7Yr
lLVYeVjxbjrW+m4Y05VT8qJ+rutnwjI9D4mvkcu/Vh8TdrO4bY3+av1qH7OMAZc7q+JSahzu7wwy
bs8f6E0+NrGsoq0C7JMkZ8lM/I2ZSkx+DutMirMPfIswxPINtARUCJtKZ9f8R9jAW5uCalBbKTKM
UwfkX9S/0lqB2atL4y5sbnwugfOBeUH8RaMbHy5go1I5EW9DN6OVEsbD9X/wc8AkbvHv9XU+SQp1
v0w8vjU7SrRm7T9FCnhIICTvTnODrKyEOCnnVXpCZ+jLp4o8qOZtGDaUmAsc0C6tH0ReoEqOZZ0+
QiPDUdSgG+AL0lXmyCB2Lp8nAiBGzn6T1gDQNPlN/nGMydNORvJZP3Q/crePEqaFAo7byho7dnqF
cuYevwQjrJMrKWoYav9Ei/was7BRjTdYC0A0ZybPwJ1TM4T3Yn+4HWcEF16k3yR3LzL0MRzpgqsW
fgiTwY2BJwOBKHhaEG7yuiS7OnJ4GEdODZYRLjBm0EDQdCQDoNQW23ScJqDVb/GQ337cylgkoMIi
t1ga8ORR2OoDpNllBCXJXGbRSQM+/MxntX9ApRrCMPYOgDdNqsBMYjlPo/JYHICDeuABNPuogh7X
Nm3JlJA07FHYmKP8rWkpDUjQIqO8sHnVdfNF0EehyCLhmbekLY6mwP0WDLOJJwZBCYto7inCzvOG
AFIB1H3JwNZ0zEp99FtOqfMZm4tGxsT4cyDTn6/aq/y3ibs3DQN+ZwshMqqXn53eC3Wsvgs7dsng
AZ6g8rnfE0Ct7y6eE4qr4JbC5e+wTrEZExoj3ttOvFDka/8NozC8XIk0Hv3Q32bZ88iUhbATPvmb
uH7kGCaBRUL1uSjlymgGQdMuCYZg3ryIWXr4opivO2SGUXbreKyCKqlcc0G4gYFAbUm8O4ipLkeR
p1sL964fE52NRDILLPTasrSZgEdwLymmtiHLvjOZh0WgiZ34S3yPmbZSbiTdJe29ogxndVlcHTqC
ojXZJGnW3dlYnb7WagvLt5umbIbCpHIiorl6t4qqam5v5GiUbe6bNQrNWhGcTbolnK1J5aAs4xKo
kpE/fRaDd4aqVYS4sb9wSuVa2dWHhTSZczWQUD0jowhw9QWefUrggXu1iLqnb/gmpB+FprfT7thJ
YFqB/DS0fpnEByiWxaeL621GSufZWTRM/yeFf8aqOy3pH1pR9F+e8OvyRWf0myME+o8AOUQk0ZJ7
zpPziB2yNK2wU6KBoS3WxT+AIqbMzim0VRegkcdndbsiYKnDyj+6Nky4dzvrxbrNtgHxOw4GbaU/
99EGcidMDeCJwlgTHShALD5FHFFv182jymBgyMO1nwo2oBEr/6HTi2nNtu223PncJCFnn8D2KQ3k
V5dV1E20dOH/mndhhwyEW3ssMKd62qCtO2ar0ruW1NP33Ghaefx7+B8YCMLcOQ9zvWlejd8Hqk4T
XwHdAs/IcCjsfDXwW4n108PHKonjTiljzL+/RqTsQ5qtqCG2dyAA2LJancJBrqi/9HnbimkyHFWB
WpY2shS7PYgKD3U7VC2JkEqxkfo9j+e+XWh1UW3uxoXrvhPBFXmBwesSTytW4I5Q5XlAcLz0oMct
mt136pwhYRwAAcg2yeA+v9J4O1Y+vZJmYiRKOTs3F/pfyJqToxCLhjny6zng4lY1XtmpdfLubGDh
m/Tf5NHK1C7sjoNi5VrYwGDvfVDre3l2hPprXRKee7/qYkWEyrrQgv+B3Z0xKL4i2AafZuTCRZkJ
lymZkXWqvIAOcwrq9piPLInwNDXEmY3+o5azr222tk/i8FZUeBYa9HBHJOaDYEZ6LgSJ40uAnRXI
UKPX/E+nvDPO/EJIhfWVaF1J/p51iV0U3Genye/r/YGHzrcKXsEVnLlQb0AMUN91/pEbsuJmqL/6
jOgdvWmd0Sh6TgPoAQWsMJ9clWhQEOLAwYN59M8p4PBy46fHVNnyyUUY/0F2liIWAFkRXucdR4Yk
Jv5RZqnRRL3dMcxidTbVinNQtodpUmFc0zUy8OA/eRJofl+IUDpppN6X4WaRP+rwHXLWBhX7QxxC
CsJ3L7dROGjfzF8G8O1ZfeL8bHGNGDWtdbICZgi5TMNJQlX3aLeHfi2St/NE14fBZL1S/k4U7GaB
WaV3xUx0skvhiKwr6I8dEwJPHFT0CsgUjgoRXGYE+mueY+t+hWoTRf5OX0aDnwWfiGFD94kPl9HX
HxjAEhOJRe1vGpq61eRq4irDw3N0M+TlVuRApERYll9b00jXKFkuPvYL0m1xXEoaz+FSh82pHdaY
ODeM2ht6CPjEqjOuPNi4tlcXtS5+LT1mSzQw6E7Cc0wZzPw7aX+QNn9WEwrdyXW0EnOhzvFhCzDk
jKeVx4AWKqC7P5NNlSvx8Jtyx1mMowvuFS7gwwAu8TeRK4JU6P/GaV9HKr9YZo5gtRfL5+LTO5JR
GB171E5Yjb3AFECeh0LGRAiSgoJvEgbKXdyjzAqaDT1y9+f1OkGrSdsrTxDHQvEjn+L1NPdUMeUC
VlVu9AMjh91WENnNVYhcUah6+lmv+IxVMgmL2iKjdqwFq5gPqTqJSRP1VO+Y8LlV9lEk+gQWbqpv
jmL1OvVqLN4PVdw6NdWwQONlg/Z8iyWylzalw2ud7UHW7R/ZelMTf072Rp3rnEhpqfIJMSytUiQL
HDlDyqNmUHXFr91SATDQoXdyprf73zuI8uRQAx1SzEMrSTTk12cvx70JBqQeoeTRHKzgjYKX+gBZ
waz/1C14ibt0CMfOt9+FJCwMvDSz1RO64OkBhHO+6Js01u1NFtZxERHBhnpz0g+vGkp0IDX62gwa
8vSj6TJn7aKLOKfPy5bow1IV5xfDPNeR55UW+ZbKe9vM2+6mzuepOGOPlWND9UkglJOZb5CFfEUu
VEhWfc0wjOlK7+4z9AtqN5APq90EW7GLTAMDoPWrnQNE9IxPCuUuTcqDFLiR/zbbaxu7KnqJ1/ae
/Z9IL602dE6aUb7Z/RZKtCg5oZne3TDGBL5I700lKm781eBOzqPvltqbd4TC+xgn8TiSmGEqX0v7
GLk0YWfPhNJH57Eka47p2XQyIiaR9ip1KS1r6C6n8fHuUYvIrFAZKgRJUSzwkXH2S3/4WHa84mES
e5pvIBjGucP+Wa4XXdl/sZGFNFLNBKrEQD4Grus7UH6mZE1QSUFhKY8RusGQiM7739zXWF3+d5Qz
/knTmbywlBRueeCRVY5MFgSY4WOH8hnNUKDz1Vt6hWU1o2vsGbk99U+VeiDCkA3lFDR8trnnfCLf
3p2sEJ8/QJ7fozapspwGDFfscwPAPQLgjL/KApyILiiemyUc78ag/qs4LGa+Wv6tA3mZTDlAcZh1
/JD6szYAIuRsCuZElMe1larhKwVj3fM3xGpjXJW31tIN6aM+UqeoA8XaxTZGv8cQV27DVjkgYRxg
yOBewUlg9RhhRxTK+uBXaZh5hs2vo3GDkbj0u+qEkgR2GQXbB/RO8YvcW7TPYBkQTXPY3XgtvrGr
wgnxb5Se9WtWSxkivX9txMa0T2EzbMER08Ngc+GnD3Uh2CZAMeAglCv4bQOy+/yxxy8Myej/V/xQ
uxZe25Ly8BvnYKO2QH/M8OKnkY0YmRYhyVXWM5IXwudbZ5aLkCJFEAPUo+rlAlot1VosVZnLsbEF
QVV4mINU1eu+yY3vcyer5r32bfy+zsHbeW8xYP7739EvsM7GzjstOGRNs46PP0D3hs009CtBkW/4
NZUbV3MgsFuR3PstM9h+PoxbmOAqHN0z+C0arv9RFQytLp4R6oI8u5Vjok8+BMCOnjZFmzIfr3A5
4YyECR538V/XFTnsFnRRRXQMDjraBP4I56q8raAn+noiqd+vMOSqlXnckqE9ymsdjO9fpoDb/2JX
fOFMrfdQTUhCw3d3FRFaEw8MbNCBDcmCad+vzOArADd70lF1EG9JRs0PxGdlQRstuxOubLvjcMQp
fnfD7RwxsEASwDs+KkMQK633KtxgXmvkuRKIZliZCDGQjQFxtfVUJ6HjKUPPceLOG3Cg6rhrCX+y
L+2w16ngD1TgKOgB4sYX84hcYWveEAlTYcKPifFgNQWQM+nr2Rpb0BUTGSNhs9rvcR3/dGmH9/Dd
di46R327+bgVr/VCr8soO5rqZrDJ5FBGJ/6XLFeumPqSGIOc5eUYQIvXaApJ4aMcZN7qNtO0gv6b
obcL5KqRjNyvj/MnJ0NptwA2tNMgNWy5D08J+l5oxSmQCH2or28IDxQ7ZCwgLGquh6iGKcFPDLFZ
54EiI2x7KlNQa2QaujmnOtfREVz/fEkELgQSz8NDzYbFus02EjDSRxZ9FjU92JQXrh6HhYJBffTL
QriONTrnVoPVf4c2IWwjrWBi8eJfe/wwUsq41Xs+9vtMU3tqnKRK0QSjL2anbWNw2SV9FkVk81Gf
9pcl9BUAw8BmneSYxZZMl1f9CqDj82toqbI9t2ejv25OJ5mxgHbs1R7Eu9cp+8MDLdvzxBwsG0ta
cFmHwwBiYmrSZ6XRZRGFhj5pB1ARuS326EhlVtrH6QbdcC4TcknZu6vlu09CYxbRzq0YbLJAifRg
sBWu2XMYTkvKjoPHLowyNERjuNAFsXT0OByXb6xq4sGkMg1t0Mc/vK1diSTGo0Gen4d76JxdI8Re
vWwArwLRxueV2VW7ozWIACfSpWC0fXP0eyrD4BDY0BawbbDkecRlaMDpCwXeQppkXzJrihuQiG7d
H81kDiJTxRyJ70h9FGM45yyq3YNTn4urfphk3RBO1pGtL2DKGqIBun+iwxEX761wiLX2NbEJLz3V
oe911caKzF7g3G7THhAYkeIOFLS+D548H/DDjmClphSgL+nB6ScY3Hdag6529Kk7Al8zq7EeDAjn
FvlalTcgSX2nIyoL32b7zAKekcDdhBmFVNgYmbQFZ2SCqja6j4+0ZZ6dUgNSNdcOp8bgzcckyunV
oujkI2y5Mwrm6fjoYEL+12Q6sVy2BcwHv87kEn6wANJomFrIYoLck4zCjgMMmO1O1wJLrT2BjMP5
q10nrF9kpUnQwYVV/oyxauuKFWXjmPn3YRpXwwP+PffpMcsj7ASi5/wmGqBBGjeO2zuQrz1Mefr2
BY7RCMvxkoUNpc5iwHUqCbsu3czzW/aCGGbSJrRBBHKEuJTfiiCukaOpNDGT6iVP9IdcCRDADqQF
SEh7SJmkVaxDjJDy3xCp7jCtPzqhKVk+AVaU2SWi7ungGNnLJrUiKPcMUNkHCLIwMhOgQuHlZEbk
r0aEn4PV+1zzGhFrEc9igFCfAXDMCmwCXmmMwVVP5CMs+oFFqxOO9V0Eba5zzkdjT4Pb9HigV8Rt
s+kx0W50S9eMDiA0hWyB8fd98i2sTyuoT7Naxm3nsqPdOhEoQZV/jq1yPDKZMpdZ+grtj68KhEtp
RxDjeiSEHTccLPNLFpe4gN4++/TQBkZqnjI14GcwHiMtwiBLESRUsWwHSVVMRTzeYyax2kJ4BfAc
NL2c2iNsoYoNMwq3OZjKoOofgUEsdGWjkfP1oeMJlOTNQ0AzSEXhxRKU5gSLCbmyi5+B1Az6w/uZ
oxgOpv6lBRVMkw75A/AbUg4T3f15x4XewoMDLd04TYYc2ZAhGhqhJwmMt/iVj30OploP1kVEXWpK
/s3UNtiO1dsmtUWsA+OcX3l4QWdS1a7bxTUwUql9RGXs1pcpwpp4i+XSWkUey8qAN9DKz4+8z9fC
l7XWteFeJe9TKn/Ws6ynrvVaPbUYLlT+HK1dtLhQz8zFIE7ITDrKiRRBycfhlQv0qPjfgR9i/otX
mIRSMWZ4St+Un7cSn0fUbE5VkyUyLIQYNfcBb5E8qYe+Ps8vaC0ffM9FwuTe4/HG9qZcRmt62/jN
qAjB/oBbM++D38sed2fagqLHrY93+svB9q8hJp+1mUgFS61+OV9sia4+SZViPumtXdB35QVuAY9T
W3fxI/Ol3bl5qat2LCGZzxDE84lK00XxQPAecKhNhmwxCZZhUTSkQdiw636J+fNAvpLJL1zB77dz
WWzSAgpGi179Khjn2BpLPZsxutrTM2ihe3IE8+CnD9pXOXAD2MCy6A7G+hcgISQugjww9Dnv6wV0
/7vkcq353L0MpCS7eYI7kVZlkg0LB3qY6mYZwHQocUPfsuyhOmTt8tWbSZ5LQTm+1zhpxfuRQh3e
JJl4yxU1c0hCps4Q1KVb5feUs7ByYegNL4N0wJ4O3Wl6tF0XRFoxIN9hGLqhr5EvNfOMxK92wc/4
aqERUHl5tW8l/Me3OeVZnO4HVXCD8hcV0uH0gUzWerwrurw+FwtCDqeSwsSXrZJO5Ve9r0vre9jV
hj3mGygLzz13VbU1zCguiBKFxy/UlxB4RTHKYCHjuEj/lV1vXP7YY1B8J07gLncu39e8o0maTaqa
Yt5jTsp+D5VUxYFkgn2v7A3rEy5OmkeU/LS2cioZWS6CyeoMkbew/ZhD/7WrQQdQye5oD9VnTPny
pm2GMcD1A2tM0TDE3RYgSoBfq3ZpoFgDaBGwAvmyJQOVgTYginG+72piTo09dcTdubl/eyLs+GsI
Spbrx9Jy70dM76f2q3liZ+st6kwYPd/mIN3axEe/87lq0jHB0XkTlGQTcJTcbRuK6nz4IizPMhCP
+DAbmDqe0EtxfbdnmINdboq/W0nWMVmFK900Dj33hC3fPDFlznUwjPyggiDodgSpm4adI3a2f0uP
FauUUowmP+42KlE5LhxFfD1OOuXpKavURy7h/n0nHBB9rm42VvEMSsYevD9w3k9dn0it79EXVFQH
kUYV9gg303W/Hn7yKWktku9i9F3S9k2Pw7i7BIGS70KmGrO7B60EnzqwC4uA/CwE5nB2jAovZ5X1
Y5/Wo5ia/NdBSZgxuDL/Xtl4xv0PQlSD2W72/WO5PQQNDNBjNIKKdiSl3GVQJ/06A6IvCQYvp7DZ
2yVgp3cQWmgKUE6i/VBwaHdUya3o52Ncyy/mPnggk+u2qrO+37+t6HuLfe7NcRwraJY+FE5qZ6Fz
IW1R9FpfSZWixvDActqF5KZnwFBWFa2KbBSYokXx+slnJWqMyKb5hM5zYTGRkzmpZfJ76zxeYepq
ZMjex1gkLyi+jZ8qx5A3h6Pr+MO/bWhQFnHhmzsqP7Ok135Wzw0HBtoR3ETwxiKuB1SnnFvCLmKh
tZuXamCbaJ42Qpl8kUaX7Va0ZvBQ1wNq9BbjDFHOxFduABU8VJfWk5B1aSVHTUZrGLc8yQuDjGPV
jEskMJAfAIJJAPnuAF4BmPOspI56At1H2G8+VNhNaxNVfXUVdQ+Zd0RrV2rUX1NgxnNVa7lrZps8
YpbwUfYTPzX5XF37juA/yFW8ASvYp/+DuUIuv4bfnwB4NN0rQpeJKz8bs6vfF/yWJ6GO03+pE7y1
nA1IrjzyZ9uC1V5FgRXt0gMZXDhPDbw+l0qMK+waIjUUhMZ0x60WZZhSTTmRuCEYY4lJc3jU1V1c
TOIvHCnF8ibHfi9bsIu+iG1tdJGErJEd3gzX4ACngjOolCVkbjiyoMTU01zqAyi074br2fjuzVPi
LL5wWJZ7r1TD78QZWjudH6bIJmiyArPT/LR4WDu6aEmdIzsjdEnvDd+nUW47voxaCYZQaJvUmWe7
jART8FYrh5zAJxhTHcMxRDtpJVEhrdbnHUD3Yj1W5Mm3xDJ1jPQT7d+0vpq4fXJXlYA2OArYtdSo
hRnBcdOXfue2jWYgedbhu6bdJ+kKT4gy6B3QJW2hDTXCMJcQq7jOjomjPQJVif+EsTmwev8UKsdE
h+4n8w2MoVgtwuZCWdaaV/lGAGjMOcWoHo/PNdLMYhYiDckGMLRLD6mFhdYmxyQm1MAiS2y8gFf4
HECbL4sJNzVb08k9DrESyGdEPcJz7Mb05wVYTvTMl80KnvOeVgmWTrSU1cLqCxYRnzdE/k5BTG+w
UBWfzmBjGQpmNHZAjeumLz/yUKbSpNjnnQB9UHeat9+4LdSt/9aozwGf7JTP1BFaT+9SprbU3SjB
o+N4hRp2W0inzQz+WiDm9In+Aspwa9MTvoqAjaeBdJutKjXnFE0LsHH9pg2Hw0/Tgi9yVjtEfhqI
K1SEtCSwfcGXTK0JwYzJuNN6UODDJFQTGZgYVOp9p9mkAXbF1SyNRDldPGmNV79JJ0bhISioV93w
w53Ve/sDdENgHL+SnUfiSA6ULr4gxAWFKiXrnfEpZpEDpbo3Gnd7Y5p2ISVCz+tiLeTkE5MSszdG
9rxY0fR676xSEScv5NpdYbI2Se0nKdkuw7KwH/dFqvRGEhNqQ+7eTVi6aQqXLoj+MzTTT9TBIfW5
fFONdZ9iNax55nd6dOKLjjTSuzN837Qp3XknmCtouaSeYz/gYnALMYvGR8adsJOkuy1Gw6V7WOyC
r+Z0BmWEyhp+tsLTIV8dsJfuIGamNNowjSTUiVOAE7dLE5YJ9LqiVl0vnGpd/TlW0L6WOzvk2FfI
VyYCuVlqfceEuCeZBct37+ZRoWG8MJxqa9N4nk53bsPEXiSS/qll86Gs9kWYdB0wWUbHZVdpmILb
HI2og4U9T4yjcawpEzvXrZE5hwkHpeWN/HJEV5PuG2NhXPcrc3Ad5CzSJjAtMvNexrjPmtMndnMk
8eF2HHuYWBd39BWwQpDpAbl4ybtb/LjoIHdR5WathOAPw/C4RMJMYPVZxhg6qpPydfui6r9ijQAr
UWpxMmAarP4hyn6LUmGBqGhMsv01npy/5pyv1Ng9LA5bn7wtgv2kH+nncOco0d5XZ17tx36elaUR
pMcWNfhGEP8yF7k0MWgBWrY1weRX0AcgW7wLiwc1CdVVeywREvHqTKD8BVuJHQPji5XjDJifrTEo
dCRHjRJB5r7QZYxRFd+DQAZWNT29KKGnEwX3HEdw/LXN3eGz6rOtZvL9/pYecJO4/C4dbCkLn5KB
cAdGNRaijqPrOCJTsM8j+NfwLMYZ49MqRNAQqSSIfhoJtVsowuj5myET728Rjpw7rrrdFLs9ceg4
7YZMGFK4bwDrRCIwVOdzP/JGPBI0f1Xm7DRjy6PFRcTUnpkA98t0Sv6QpYiGTottI9+u263P75xk
QxobRG7ayBy5kmZYJUg/UFduMdzIEkx+mYuj/owSIn7SSZDXU0xHCsTyncTQMfclubzxyhe4YU99
6awheA7xGm4smr2d9zB3QDHPy0298bscD1zmxbg2qUm216+j2qtc5/3I4kBPCTTXfyjGXFfnGJqF
C47azELdXMgaFbhMj0gt1K5jAMCBZf3FPLc3REzhplVHhUQOeMavh6TIILLlge2ppX/t4U6DsEnM
gnAYXdysgB7/0GKMEV2YV1ZCoX6378xozpFQkM21WGcOnyvg1g/1FP4gf04MJcWQa8n2laiwX1FV
uhYVS9meqp5yc1VennOOAkZTKNf+54Ys31sc9bRpy192viAxPAuJ8Wy6wmuVVO6UmPLOSUDgJHgY
xqmeJxm2PHttZoYjHAUOVR9M2fMKoiHcYur2NoPCqiX7qR0K5kscVKNF2ZdUixOrUjg07t4g4F5A
E48kODYauqZEOH70wWcTvXEaZSbJb4y/b7ai5/oFQMJqeT9FEpdMWXYCi+pb+mv+wfDUE/3UaItl
xLMeB/REqe+e6p3ZY06IOINfs+R1vOq7mAkh57opVu8nWE8nYC5CDP7f3Bm/rNYcyYvXzPiFDCJO
Ay5s9oMIRb6sE2jE0GNEw9+smNPotED5T5/+Jej+qECDxMx0rLILNQazCyZ/6/jyeeP3TgYp2KiM
CovRB66I2ekuWj70kef9uJbOFT53qHY83GdBAXQcUFBBDmSNfDH/6M/8ql9QzIzwfC5wvmK3/XtW
wBD1zomwI0UeNGtAUyI3TqybJxxDpJR5/82xf2a4jcwRBV+JWEN1LCsjjFyMTGTaaFZKXL4iSPd3
+opFzA81IugMpcp+OoI4uk5q0vszms1IVVauoSIiSegi2upkggBqSA/L7ZDxG84xLwUzxjecXidv
J9f7xzUlcjGV+WbzmVSFraerPTz6V4YFgau0Fen9/5P3tYhrPxGg/HdOIQCtm+GtRNli9J9W2bLj
9m0gKeDLn2IKyd0YZNM0HRTNXH7GR0oRi1DnF254e1Jw6bHLuqss54CG94tb3Lj9wQ4Ze2VvsjKL
NFX1rClSfsXUpT3csP/Qmop4IYVuHjA1rA5Fi4sRsW+0hb8WSu7k9EHCDgEH5L8XuxL0SOYXpfXH
84KXom9dlQg2flEvpxDG29zQxXx1O+RE6glzOq/3PtQdG8la8aaaoEkRM/qDPFhccFSCAV1QHUyS
mX76uKDwtzo+I/tnKYfnaamxqZ22ohWyF3gbIrDwOh+7/vLl4Nu6GejaCDGK3y8KO9+qKiucQe35
qSTjBQBqiKTlNOu/PrQFSZHBIG42e1BaE9+2CHvO0Eqi3+8h1LASqv2UMnXFQ6Yml5sbXaivanMO
kCwTLYgB0Bt6dMZ4wrzVCVonn9+ueloG18rc5E9/nIBmG+3rfEAZM4vJOk9/imNcCwG9k8U/QJVh
c1GeajSQc8dDsI6mL9ZW+N8iJUbJU9acPwFHEeoQYgbd61c5hgiftFlD41iaIX00T+qbiwfhzcX6
GJg3OzgSpUMMBGryw4USaNIJef4uhgW8eK38pXlOUmvopnG2juPh0YVXYcxPqsYHR3SyEA7AipZA
A4w2ZYRMDua9KwjXas3T2r048QRVOmdf4wgxkHwUVbocBvlEvDG5fJAyawh8UZpq5G0vJbeJuDVI
S7ZbbIq/hCpGtZzklr/70zm6LFRwNNhyPAUqE8oWju2JaNakD+5Pn5wxzR/taT7hxHiPqdrouMXW
E7PWGsgmtdiygoXx2/ibEWVN1Gh7cYqf4/7cbqXCtEPeBIvrLjsciKNj58m+tbngkiKS9P0oVJtj
HLkOI4PSwDsGBWJpT6yAV/SFBHUdrfaQXu4KfIXl8rsVFbRXfsFGh+/TU0LcEKUKXd0SR3eNTCht
9/MlIUk5UOfbnIbyIBL4II4XysxKkfkzump/AmwNLUIXI9kn398KteRDaJyc6+Pp69qpUllMnqT6
NK12hhSyfm/m0JIqSDmOk3hCqg62AQUR3xHo+/fqwof37UMyKbzXBZo0FbYZTZcVgTAxQTwqIoXK
awXEWGUXYxvi7YTw5/KSzhxLFnV0gZ9OMcx/xgQKZNPc+YnJgwDl4MLpiu8LElX+VqgsAPO7n5nt
H7DfTXoUGnfFfOea41qjg1oBQU69HWuxHIe4o8MRyD7wjxcQSaroL88oYaS1d3dqKlBlp/zGVEFl
wG8AK9YAJkRgPNJzQJ3l6qPcfggJ0WM/UVNH1zfvD0MjFCS/UnVSa13atJFNTfD0HEub0ANd0mSu
DSE95/KT3FM9ahucQ77hngtDXdZ/Ug8NDU+A67CZ0uHcAPIMEda1LWj9ZDkh3XQt8rCHQw8mmSAh
1QRQhq2rapqMsT4HWZh+UVIyzvAMx7JDS2EZS1ZRYoHC/n9eaTk921JTVWD9pQtOf9ObrX5Qyhtv
4rLwPUAJCVpPt/QiDen6AmYiMhYXCP2Jhffljyznxhg7UI7OdNzO2zvVtgEX0QHlgdy/4y2QETac
BI7vjFS6B9IwzHgjkZAnDfwpghQnbhQYHa7/cHgMvDwEu71EUnIcDN+zySnegsH4izF9sykOM86K
ljIZiLYAwLbRgDkwa52e2ih8tgtsv10PpdzBG/5q216k/gdQwh+UmJX87YgR9E4UtN7R4l22/lwl
yGNH7c7mv+kOLjICibZ4+nx1KDEYjav8iG/haqe5q88bIedhaSShO4lxyvxuuGDw3HOpEDR+ccDR
1saWssil0mRMK0FvKVv0XNshAHiD66+5CfY4i+prv3MFlBj7Yw8rkxKCMvgAfRJEk3vuwxcXPE90
OwFrQCt9p3fi1sEduvdgdaRjEi8+vbYYUddk31ykye47rg2Vv3b7Ukuqg7Kb/N7iz6SaBY6UMRmV
iDJAqLv1jXGWtqwMtbfbzO1Fbk9z51jPSfl6s/kJEriEeMz8pTKKuAcy1qmLox99gEHv32uLnXK2
3LHjX3VZvv6crbZMd6o5uaxaFCgoo9sh0UXNcQMz+obXeJCjJ5zS6dbFFtKHvl3X7HYnOGsL7h50
/b5ZspwFrAby+zCwg/Ko6W1Aq+a4+HGDCX1HmdhniDyMCdpZhCidD/qGJflaYmPeWIZkpU4wrgPR
nKRqq8j2kCtAi8oCWfqM1Zp/vc6WpimVzYXiGCf/6t+n6DBOzMgOBMH5U/GgFDpGbyPUDOu55I1Q
GLd5zH+qZPPWnV9x6rRLTFjxw3LnPA6DMRzEQqme217lER/RE3LLwL3e9eeySZMr1Xgn41yLgnkz
dQYUuZgT6q3kfLFeJ0pNCMrX4Z24kJ+xxYQRglb+yAxDziXT3R/e0Zc1E9+0iY917Qja6Ea14vr/
1ELkYU3eoYGPnMoEq7klfFE8htvdneEAiV9IAUAY3pv8lxTTNXBr9Qqni4oQlt6ecR/JpST1AuiY
x7DFkrIlVKz3UK30nm44whXSv9MJjzxQPCQ1OXW4bd5TALLrKurHSR51QvBtxR5JwYZLICo1ZRJ6
rZPG8ylmRMYnSCxApfWp31P2KapvVHMCCTGAKMW5KQITBrQ9qWcLwvGrIR8/A99gly/KlvzKjt89
GEbxWi6OjW3HOSacGL2efSY7FgIVYYOWqbvm864FzdF+toRpkaL6e74WBsAcb6g5VoYqljXrEb9M
oxZEXzeuW5RGuqSdWg9WxvC2RMBbtz3WJvLQGMug7llv0Np9MDacLTEH4HF9zS149J5MF2u/ztQb
4uLwG8YOl1Ljo997gfuzt6ZnyAvzlNW+8meE/y2nz7ElXr4JLwUvC+G9xu7FOtSm/Zte2MAj7UTS
s0q9LMRODeIShUsWwEDTl9O0eVRf8DLCE2mdfAuQFUW5Gp8KPboAhEF65dlwVyb5EgWuBGm04tP4
adyzCi2Se/jSVJcNrMlz769XMhE2GTO5PI8XPBZc44iVSeNdik5reB29yTHQ7wEjjTwEGO2bKaI0
T5fDH5dcCqeOc+4mx3grvvNL5Eg4dtHaUfcnEdbK5YXz3v6rMfEvxXRoCcOPHokR6EazygpkTDT/
57ymveZK5yU7DFl8QierNpzQsAPCREipC0HAW0qPudMhOXGi+4yG1L5AknzslMW6RJOyBmiPbhwr
pav0bi+6Sj6YImqh8UUiI/xHKb9KlK42YWVc8xeCLPWxiob8KGXBXfW6ZYT5uthDO3V+A5hgNRgg
4XbwgZRbfEozTU28skb6zskasU70pB436j59aqloRgkqc4GHUZiPz2Pz6ikOQwQR1pWSs7y3GQo9
iBLGoiM8OP61xbUHRc1NVGk+Zum4Gyt5rEpOC8Kcub9ECneCYIjJPqVYviV6ohg8VsNBkFvcOkeR
TIk0LjbI8V7MYPYCACEWaJqrXS61gyhFiQBrfEyBBQa58ij1NtxtDWqpAO/EDtramLnlfBVzs/6V
9TxkI9//h8BVW0gNpJpvXGwjcdggc50s6LNNO9iBo0JgNVZpzZmKZonRi8GHnQE5v5lwR33ID9Ey
ZdCsnIL7DbvY0PF50ovi9BN/4z+zE1XHvK/Z/fTjLRFZQuyV5EZmbnHpXlcrtDEfmSvbolsSxMj2
0qVhpIDyMP6x4gqxmdt5VSHFLRJRV8s5dyMsjKxzc4BVc2JXor+Rf+nEabZxB5msbXLlQoxBD6xI
bB3QJ351FIyh1Gqj7U14FRT1Y+oXxRdtDC+eIpJDUwG7pqCeZ9yYyabCdeOz6HcUWTIhgkbEQ2ST
EHjCVfkF519qJ39AmJiYVVhe1CwypzaIKhiZ4XSS5kolVSIJ4W2IhXERbEukXR0jnURvUXCMlBNg
KaReLdFEQzcmuNC25/7yNRLviV2rE5MzvVpmagHhBu7Hi4nvRpameHjXeWubsLnpElLwKaK33sCL
vatI7/uqfWhH3ajLVfAG0JQN3/6mKP2OqZVQMffiyBriZdfYLABwLPIjQv178iao7NBSx2Nw0oou
MGymxmu/tGg+Ox6ralrzqDh1NfPA+pbrXV+EIFwxR/mPhtEvEaDGmzEk1gjFv8uMSszzE8H5vrcl
o80eRNcq5Ur4OyUxc/n4SwPJ2gpGSB9MkdYx3LFqmOtvsT7CTTYO9ZRvQi0c+fjV5kjg7rz7Xp3w
2BprgMVBoyoYtjLrruleac2mm4o0t4Q+Jr3BILMwNYzJS8bJHjxHbgaJhfLTwmpsuuij3FtidVH3
yRiJ7ee0yeOX1xDGQ7LFK+WbbdIXz+vTI7EjdFFWll7qqvM+rxRRSCButsGO6EWvv9P6SM1JMiJS
7pvBY6Kg4x1Rdqc4UY7ARcCNF+3wnUPkTebmaiTnq5JsDNIJZUbrrdjVO4k7fUXQFZNv/JBl6nKz
WqIrW8FSjjOFIbVjiIa+Vfd/B/aFZgPLNq065QGGL4lWmrymsjVV9GOEoPAH4Wv6t/k7/VFRpq6C
pVh192gezB0/RAVmNiquPsI/0g6b8/5fSr/E2VPvkKWZj/AVOqxjFNiP92G3De+YMRKZOGgQuNNd
qgFn/Lgzzzl46l9HFHLfuRBnTdimT4XSBs/7iypIHvtejEzmYxQCdtHgbOk9UouyOVZmrn1tpY9o
H7jQvNM6Ikf8SktckubuT5Z1WBOm+piMhiLIeHzdH+/o0kZohzoq6RMyszxcwJ4MokA2fXn+lDJq
F0Rv814fNeyN9foVAfl9W9t2LdA3BnU8Nib7+nx+GYV9A3wwQAyV5WOfDLV2F59EAlWEY82HzFFK
cauCVSSu0e6X+4XaGK8vDaiaSYEdvfZTh3IdTTKomIiiMFXn9t3AtVK7uGucXTVLWfzMYTrqqmRB
mjPpW+7jfBGgnarAObDtsZAygf50nqvoQ1Bc/AmFvphgyZPhcnj36n5vK5pz9Oy4CYA7tvGuYIjP
+vYXY4vx1QxxYwd/WT7S55SWixz6clWq/neiZoq+WnE8smrbcLBUHvGVbgi1rTaclC60bvKFCSC+
FAHXbzTJ3L+8OPmbLGq/jMkpymgZP19su7QYifzq/UxteekNSZ+7qn35J/W+uzrQKgNjs1Fabwp7
IPco/J/NgGEL6rv6YtCyWzzLFVTr2F1ZXonPMwB9exIC172kmZqAQurZt42N8fsli0VQAfbHo+zU
VwYoy19tzYMlr/NHSZkzc5J4isUpk8GRIOpBu4QdJ4huOFGGl+nMtIBrPqH91iSKzt2oqk4Pjjqw
WEWUoGIZ5dZzpzhEolkDycCY71r0PbdCmFON55Ko7BLkgUx4Mh5xyxUbNCpLVtJG2XdWPuRBVGX5
yPfHG7SoPO4HQTlC2TkoYva6oeZfA1StRx5I+gmA1kh78ZLnFT9qz+D6DgsV4EdNcWQsTZS3MTQ2
8zydcaOoahhvoaRFTZPWWa7Rs2oaz6uVNMSYfvBMO05ZQTAMB2dnKCjOwTMyiXxB6ImNFaEL2f3m
m36Nd040h9AlaL47qxrRdSctb2nmT7Yo4SYg/v+w+/8OfcFDMOfGvm9MqpbDyUoSza2BrxA8QHLZ
FVVfztJsseIPqdcMhhGoAk9GTq5bpJSe2TqqrXQ4deoP3y4iA0WYtMM24ijUOx3N5Q/8FC3nOHVk
XJWXBcQsbmCIiN8jTCtQH+S2E5dqRJN7Z8pgGSMIq8NcDqDiK/sJmppHIeAfz2MwiM84MFRIUHD9
53abTQhbk59aI3LrpHjGQnKIjvi63euL8/sOuYi++14IWpMSPWJLdczv9IE6EOJs4lzXagpLN17q
xLL6ca986WwAWnay7dh3SehbsjwJjc0pUj2xZaE0XMLD5HQXRtDcqPC85p531z0PjIIZCq9sEjj+
zJDiPUPSWu/9jtsrEb0qAQN//CVGG0vgsU1BBSt3U2GABZLneqjQUVV0PzztBYGsN486uVZlpc3c
1PiHE9B++RVfkxwLLAWLR62dBHSbwn6G9Jcs07gu93CphU8tf9wJ12G8Gth2ek1riPFOvlX+BNu1
6PHB5HMS4XH++Qds8IOCH2VQr1mODALktTYVJwnoCi8dAezxSgUC0/LLIE00D2fq84y4sYsZiVwL
YcfXQUb7+agR1+7ppb3X8vNIHzEhE/hD8y6yhaX2a3kvtsh5ZoP4uFs2sKGQHE/fvXc2270h+arT
t8NBYgN6sAo3KYxn91nS1XD5FlWsWfKSY2V5VtwV5I5XKWsjpk8XXZNzar4dBVnpju7cA/GIR+1B
dnJ1xI939Md09uE5d1NA0oQPYYmKmeN5bpoFgUNzziPTi0Fn9RT7yu783WC+5q9q+rSQRxJe6ycy
6N+hjB5JAoELB+pFpOZaqH4FTAZyUmN2EHA3+dtJg8QtOwaedR4K+yV/D7rVSEh3kTsg2Tpcq0AQ
pfjfNKSpU7EM5jH0YXIOwOycp2DRw+wYeNdA/awFbz82Zlc5H3Dhds5sm0OWXcVSHGOJFottNKGY
wOpke1//3OTd28mll+1vJeipxpc1ikB3cNTgAhliRW8AKl1gzsYJ6fOjUeTVNCmOGaOqMW9hFKGu
idDoqg7Fe8WEhUM0E803ZZVoOCkNignYxH8mdpSh5xSosTNjJi0jWwHI5sx06XQSt5vgQ3okFi4a
/aUEAPUQWvtgnimUGeC5vMrF7tAXw0vNU/TFN0USuRQYYjG5WrNJgiZGg7IPuHA9F144fd55cXV1
9/Hq2U1ebV5wbELL2afgJNPf9wuHLLdyNO7AFc+/BnqRbW/h9Hzff8GUPPRJmQxQcVA1CdxGEFiO
M+y8NGSoUARfoTPk5JRJviPXdaVBNcwIg5NNfgJDXTUbkVexlmUeWs2OIaAbidJNWeTM+87m7lxm
96A20QFFXZuIhiYC7tQXr8Cyov9XSREVOTAYEwwyqVeibWRapU6J9puOSfTipiH6XvnlYyjB8QjM
6mgjxeipNUfig5vyee8ijvi5jsW1lYqs/yoRz6v98h5M1iYEmBtNVUEevySft/bRCTpU8vS5iO4j
PJVAqkMIoZP2YwsxJqJXmqL7XUfnPY0x7eMMfUCWcgTrrjzyNh22aNrRBpYSJr8EncsBHY/kN7/i
oD09nplhVfkvKt+oXrXpoQTiYLsI130YqKhKh8+5/7YAg4j86U+KFhS39ieSapQhrAOlZ3ZFdHIh
S3wAOs35NcuyXsY2bcw58P4wBiIQ/GYjsVKXRf+SliWoPoHracYIrIs3BTISeZk14zrCPALmt0t4
qWFhNc2rVi4EU4zXUWXQpgPop+wwcCbeGKNR/hWHHjilPtbLf5NssE09f6YUuWt1LO9vQobVDJIS
ZTNw2eV2ncX+rqAJ9rxY/o+FX2PoGvAXhaAveDMd37+sNlN2SXA709TLrYW81Ne7P53QOAjhspwI
gGY2hGq8pcGSufbnQJw2obR1mtxld6hupl8wVmfjAnguYMYHgZJhxzF7jiVbuyV73vNiyqhxtYt4
lQRumpaCxIIyAcL7WpcOTVMZMfRGFawxlIJ4uwE40bAt/A4158ok3e/7cz4YtrDGGm/jr0cPCEzG
gaUZAUP6XcW6MamOAZiAK8cfLlhUdZ0TeJICLuPhcgijBL4Pv8teL+27K74hOyL1XSyvDzypzx1m
MPdS9rFHlDjfqdacIAXcAN8eSAyRk0DGK3092LrGuR/jm8IliQjQ0fXwJtwmtWOe6cv9BEvRlVZP
OEtBfeXEEeNmnrZVq5I0AvLGR41Yl+zgNm36DQUF4l3ME89G1ZtHFCy5UjAlhVT4C82Lc45rtEhF
kKng6+/hBj7wC2a8/Z9HFmC2kU8mkm4EFIVZetnixCktieCoVXiEOgzBAyj5WNqh7JruOIBStVIa
JuCRCwTvFcPDwZIHbknG+6RfFTEjOpHyGNlxsKJCF5/GSIUEACEGDgV7m4syCYCjWgVopmw2SvJn
zzmLAmLhfEXtq0CQkhEnuhgoKunKTnvvkv8PhZ4GbaV8GG/yajfXEmHBWQ4hHjrp6Aywq3mOKw0z
mxRIxKCi4VttmqcLS8Eo19wgmzSUqU7dFs3gyx/FRyoe+FW/+i5eZND6C3H1/IeofMPkLgT5sNis
Xsr3fDROdiCMpe6s7bWgq6paVXum7uw3nWjifXfLFc69zr8Sru+3VBHA6k9CrOzRNmR8x4jKUDSN
JC1rKmatb7thMMFKPjqPN5RA8Nb/3I/knG94bNms7ywLiiClATi/QcgJXp8s6V4rdjx96zCu3oOH
RmiATpvYYmFS3WPcB/YWzo24oEEYYih7IfsJdYzyYk4id72rei6qJ3nSqVfguuQwTXJ+1TCGWcO/
xgQs2JVMVnojbBoJNlCBH6WKhH6PlXpPggtN4tU3a8chE79xo3M1odQeY8Ztcp82yjHGTFIO6JD2
qSHfcXAb2hA0ZG7T6eN5/0kn8CQEiC2gyGPicP+19TNh
`protect end_protected
